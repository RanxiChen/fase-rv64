module Queue(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  wrap = enq_ptr_value == 3'h4; // @[Counter.scala 74:24]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 78:24]
  wire  wrap_1 = deq_ptr_value == 3'h4; // @[Counter.scala 74:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 78:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_io_deq_bits_MPORT_data = ram_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_1[1:0] :
    ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      if (wrap) begin // @[Counter.scala 88:20]
        enq_ptr_value <= 3'h0; // @[Counter.scala 88:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      if (wrap_1) begin // @[Counter.scala 88:20]
        deq_ptr_value <= 3'h0; // @[Counter.scala 88:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NulCPUCtrlMP(
  input         clock,
  input         reset,
  input         io_cpu_0_inited,
  input  [1:0]  io_cpu_0_priv,
  output        io_cpu_0_ext_itr,
  output        io_cpu_0_stop_fetch,
  output        io_cpu_0_regacc_rd,
  output        io_cpu_0_regacc_wt,
  output [4:0]  io_cpu_0_regacc_idx,
  output [63:0] io_cpu_0_regacc_wdata,
  input  [63:0] io_cpu_0_regacc_rdata,
  input         io_cpu_0_regacc_busy,
  output        io_cpu_0_inst64,
  output [31:0] io_cpu_0_inst64_raw,
  output        io_cpu_0_inst64_nowait,
  input         io_cpu_0_inst64_ready,
  output        io_cpu_0_inst64_flush,
  input         io_cpu_0_inst64_busy,
  input         io_cpu_1_inited,
  input  [1:0]  io_cpu_1_priv,
  output        io_cpu_1_ext_itr,
  output        io_cpu_1_stop_fetch,
  output        io_cpu_1_regacc_rd,
  output        io_cpu_1_regacc_wt,
  output [4:0]  io_cpu_1_regacc_idx,
  output [63:0] io_cpu_1_regacc_wdata,
  input  [63:0] io_cpu_1_regacc_rdata,
  input         io_cpu_1_regacc_busy,
  output        io_cpu_1_inst64,
  output [31:0] io_cpu_1_inst64_raw,
  output        io_cpu_1_inst64_nowait,
  input         io_cpu_1_inst64_ready,
  output        io_cpu_1_inst64_flush,
  input         io_cpu_1_inst64_busy,
  input         io_cpu_2_inited,
  input  [1:0]  io_cpu_2_priv,
  output        io_cpu_2_ext_itr,
  output        io_cpu_2_stop_fetch,
  output        io_cpu_2_regacc_rd,
  output        io_cpu_2_regacc_wt,
  output [4:0]  io_cpu_2_regacc_idx,
  output [63:0] io_cpu_2_regacc_wdata,
  input  [63:0] io_cpu_2_regacc_rdata,
  input         io_cpu_2_regacc_busy,
  output        io_cpu_2_inst64,
  output [31:0] io_cpu_2_inst64_raw,
  output        io_cpu_2_inst64_nowait,
  input         io_cpu_2_inst64_ready,
  output        io_cpu_2_inst64_flush,
  input         io_cpu_2_inst64_busy,
  input         io_cpu_3_inited,
  input  [1:0]  io_cpu_3_priv,
  output        io_cpu_3_ext_itr,
  output        io_cpu_3_stop_fetch,
  output        io_cpu_3_regacc_rd,
  output        io_cpu_3_regacc_wt,
  output [4:0]  io_cpu_3_regacc_idx,
  output [63:0] io_cpu_3_regacc_wdata,
  input  [63:0] io_cpu_3_regacc_rdata,
  input         io_cpu_3_regacc_busy,
  output        io_cpu_3_inst64,
  output [31:0] io_cpu_3_inst64_raw,
  output        io_cpu_3_inst64_nowait,
  input         io_cpu_3_inst64_ready,
  output        io_cpu_3_inst64_flush,
  input         io_cpu_3_inst64_busy,
  input         io_tx_ready,
  output        io_tx_valid,
  output [7:0]  io_tx_bits,
  output        io_rx_ready,
  input         io_rx_valid,
  input  [7:0]  io_rx_bits,
  output [7:0]  io_dbg_sta,
  output [7:0]  io_state,
  output [7:0]  io_cpu_state,
  output [7:0]  io_opcode,
  output [7:0]  io_rx_data,
  output [63:0] io_buildTime,
  output [7:0]  io_uart_buf
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [127:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  wire  event_queue_clock; // @[NulCtrlMP.scala 76:29]
  wire  event_queue_reset; // @[NulCtrlMP.scala 76:29]
  wire  event_queue_io_enq_ready; // @[NulCtrlMP.scala 76:29]
  wire  event_queue_io_enq_valid; // @[NulCtrlMP.scala 76:29]
  wire [1:0] event_queue_io_enq_bits; // @[NulCtrlMP.scala 76:29]
  wire  event_queue_io_deq_ready; // @[NulCtrlMP.scala 76:29]
  wire  event_queue_io_deq_valid; // @[NulCtrlMP.scala 76:29]
  wire [1:0] event_queue_io_deq_bits; // @[NulCtrlMP.scala 76:29]
  reg [1:0] cpu_state_0; // @[NulCtrlMP.scala 41:28]
  reg [1:0] cpu_state_1; // @[NulCtrlMP.scala 41:28]
  reg [1:0] cpu_state_2; // @[NulCtrlMP.scala 41:28]
  reg [1:0] cpu_state_3; // @[NulCtrlMP.scala 41:28]
  reg [63:0] global_clk; // @[NulCtrlMP.scala 55:29]
  reg [63:0] user_clk_0; // @[NulCtrlMP.scala 56:27]
  reg [63:0] user_clk_1; // @[NulCtrlMP.scala 56:27]
  reg [63:0] user_clk_2; // @[NulCtrlMP.scala 56:27]
  reg [63:0] user_clk_3; // @[NulCtrlMP.scala 56:27]
  wire [63:0] _global_clk_T_1 = global_clk + 64'h1; // @[NulCtrlMP.scala 58:30]
  wire [63:0] _user_clk_0_T_1 = user_clk_0 + 64'h1; // @[NulCtrlMP.scala 61:40]
  wire [63:0] _user_clk_1_T_1 = user_clk_1 + 64'h1; // @[NulCtrlMP.scala 61:40]
  wire [63:0] _user_clk_2_T_1 = user_clk_2 + 64'h1; // @[NulCtrlMP.scala 61:40]
  wire [63:0] _user_clk_3_T_1 = user_clk_3 + 64'h1; // @[NulCtrlMP.scala 61:40]
  reg  cpu_raised_itr_0; // @[NulCtrlMP.scala 65:33]
  reg  cpu_raised_itr_1; // @[NulCtrlMP.scala 65:33]
  reg  cpu_raised_itr_2; // @[NulCtrlMP.scala 65:33]
  reg  cpu_raised_itr_3; // @[NulCtrlMP.scala 65:33]
  reg [1:0] last_priv_0; // @[NulCtrlMP.scala 66:28]
  reg [1:0] last_priv_1; // @[NulCtrlMP.scala 66:28]
  reg [1:0] last_priv_2; // @[NulCtrlMP.scala 66:28]
  reg [1:0] last_priv_3; // @[NulCtrlMP.scala 66:28]
  wire  _T_6 = last_priv_0 == 2'h0 & io_cpu_0_priv != 2'h0; // @[NulCtrlMP.scala 69:37]
  wire  _GEN_4 = last_priv_0 == 2'h0 & io_cpu_0_priv != 2'h0 & cpu_state_0 == 2'h3 | cpu_raised_itr_0; // @[NulCtrlMP.scala 69:97 70:31 65:33]
  wire [1:0] _GEN_5 = last_priv_0 == 2'h0 & io_cpu_0_priv != 2'h0 & cpu_state_0 == 2'h3 ? 2'h2 : cpu_state_0; // @[NulCtrlMP.scala 69:97 71:26 41:28]
  wire  _io_cpu_0_stop_fetch_T_1 = cpu_state_0 == 2'h1; // @[NulCtrlMP.scala 73:77]
  wire  _T_11 = last_priv_1 == 2'h0 & io_cpu_1_priv != 2'h0; // @[NulCtrlMP.scala 69:37]
  wire  _GEN_6 = last_priv_1 == 2'h0 & io_cpu_1_priv != 2'h0 & cpu_state_1 == 2'h3 | cpu_raised_itr_1; // @[NulCtrlMP.scala 69:97 70:31 65:33]
  wire [1:0] _GEN_7 = last_priv_1 == 2'h0 & io_cpu_1_priv != 2'h0 & cpu_state_1 == 2'h3 ? 2'h2 : cpu_state_1; // @[NulCtrlMP.scala 69:97 71:26 41:28]
  wire  _io_cpu_1_stop_fetch_T_1 = cpu_state_1 == 2'h1; // @[NulCtrlMP.scala 73:77]
  wire  _T_16 = last_priv_2 == 2'h0 & io_cpu_2_priv != 2'h0; // @[NulCtrlMP.scala 69:37]
  wire  _GEN_8 = last_priv_2 == 2'h0 & io_cpu_2_priv != 2'h0 & cpu_state_2 == 2'h3 | cpu_raised_itr_2; // @[NulCtrlMP.scala 69:97 70:31 65:33]
  wire [1:0] _GEN_9 = last_priv_2 == 2'h0 & io_cpu_2_priv != 2'h0 & cpu_state_2 == 2'h3 ? 2'h2 : cpu_state_2; // @[NulCtrlMP.scala 69:97 71:26 41:28]
  wire  _io_cpu_2_stop_fetch_T_1 = cpu_state_2 == 2'h1; // @[NulCtrlMP.scala 73:77]
  wire  _T_21 = last_priv_3 == 2'h0 & io_cpu_3_priv != 2'h0; // @[NulCtrlMP.scala 69:37]
  wire  _GEN_10 = last_priv_3 == 2'h0 & io_cpu_3_priv != 2'h0 & cpu_state_3 == 2'h3 | cpu_raised_itr_3; // @[NulCtrlMP.scala 69:97 70:31 65:33]
  wire [1:0] _GEN_11 = last_priv_3 == 2'h0 & io_cpu_3_priv != 2'h0 & cpu_state_3 == 2'h3 ? 2'h2 : cpu_state_3; // @[NulCtrlMP.scala 69:97 71:26 41:28]
  wire  _io_cpu_3_stop_fetch_T_1 = cpu_state_3 == 2'h1; // @[NulCtrlMP.scala 73:77]
  wire  has_itr = cpu_raised_itr_0 | cpu_raised_itr_1 | cpu_raised_itr_2 | cpu_raised_itr_3; // @[NulCtrlMP.scala 77:42]
  wire [3:0] _event_idx_T = {cpu_raised_itr_3,cpu_raised_itr_2,cpu_raised_itr_1,cpu_raised_itr_0}; // @[NulCtrlMP.scala 78:52]
  wire [1:0] _event_idx_T_5 = _event_idx_T[2] ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _event_idx_T_6 = _event_idx_T[1] ? 2'h1 : _event_idx_T_5; // @[Mux.scala 47:70]
  wire [1:0] event_idx = _event_idx_T[0] ? 2'h0 : _event_idx_T_6; // @[Mux.scala 47:70]
  reg [4:0] state; // @[NulCtrlMP.scala 140:24]
  reg [9:0] trans_bytes; // @[NulCtrlMP.scala 141:30]
  reg [9:0] trans_pos; // @[NulCtrlMP.scala 142:28]
  reg [5:0] errno; // @[NulCtrlMP.scala 144:24]
  wire  inited = state != 5'h0 & state != 5'h1; // @[NulCtrlMP.scala 145:46]
  wire  errored = state == 5'h7; // @[NulCtrlMP.scala 146:26]
  wire [1:0] io_dbg_sta_hi = {inited,errored}; // @[Cat.scala 31:58]
  reg [4:0] opcode; // @[NulCtrlMP.scala 149:25]
  reg [2:0] opoff; // @[NulCtrlMP.scala 150:24]
  reg [7:0] oparg_1; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_2; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_3; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_4; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_5; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_6; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_7; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_8; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_9; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_10; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_11; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_12; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_13; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_14; // @[NulCtrlMP.scala 151:24]
  reg [7:0] oparg_15; // @[NulCtrlMP.scala 151:24]
  reg [7:0] retarg_0; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_1; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_2; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_3; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_4; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_5; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_6; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_7; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_8; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_9; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_10; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_11; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_12; // @[NulCtrlMP.scala 152:25]
  reg [7:0] retarg_13; // @[NulCtrlMP.scala 152:25]
  wire [1:0] opidx = oparg_1[1:0]; // @[NulCtrlMP.scala 153:25]
  wire  all_inited = io_cpu_0_inited & io_cpu_1_inited & io_cpu_2_inited & io_cpu_3_inited; // @[NulCtrlMP.scala 156:51]
  wire [4:0] _GEN_20 = state == 5'h0 & all_inited ? 5'h1 : state; // @[NulCtrlMP.scala 157:51 158:15 140:24]
  wire [1:0] _GEN_21 = state == 5'h0 & all_inited ? 2'h1 : _GEN_5; // @[NulCtrlMP.scala 157:51 159:49]
  wire [1:0] _GEN_22 = state == 5'h0 & all_inited ? 2'h1 : _GEN_7; // @[NulCtrlMP.scala 157:51 159:49]
  wire [1:0] _GEN_23 = state == 5'h0 & all_inited ? 2'h1 : _GEN_9; // @[NulCtrlMP.scala 157:51 159:49]
  wire [1:0] _GEN_24 = state == 5'h0 & all_inited ? 2'h1 : _GEN_11; // @[NulCtrlMP.scala 157:51 159:49]
  reg [47:0] hfutex_masks_0_0; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_0_1; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_0_2; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_0_3; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_1_0; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_1_1; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_1_2; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_1_3; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_2_0; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_2_1; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_2_2; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_2_3; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_3_0; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_3_1; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_3_2; // @[NulCtrlMP.scala 162:31]
  reg [47:0] hfutex_masks_3_3; // @[NulCtrlMP.scala 162:31]
  reg [1:0] hfutex_pos_0; // @[NulCtrlMP.scala 163:29]
  reg [1:0] hfutex_pos_1; // @[NulCtrlMP.scala 163:29]
  reg [1:0] hfutex_pos_2; // @[NulCtrlMP.scala 163:29]
  reg [1:0] hfutex_pos_3; // @[NulCtrlMP.scala 163:29]
  reg [47:0] hfutex_match_reg; // @[NulCtrlMP.scala 164:35]
  wire [47:0] hfutex_set_value = {oparg_7,oparg_6,oparg_5,oparg_4,oparg_3,oparg_2}; // @[Cat.scala 31:58]
  wire [47:0] _GEN_26 = 2'h1 == opidx ? hfutex_masks_1_0 : hfutex_masks_0_0; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_27 = 2'h2 == opidx ? hfutex_masks_2_0 : _GEN_26; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_28 = 2'h3 == opidx ? hfutex_masks_3_0 : _GEN_27; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_30 = 2'h1 == opidx ? hfutex_masks_1_1 : hfutex_masks_0_1; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_31 = 2'h2 == opidx ? hfutex_masks_2_1 : _GEN_30; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_32 = 2'h3 == opidx ? hfutex_masks_3_1 : _GEN_31; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_34 = 2'h1 == opidx ? hfutex_masks_1_2 : hfutex_masks_0_2; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_35 = 2'h2 == opidx ? hfutex_masks_2_2 : _GEN_34; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_36 = 2'h3 == opidx ? hfutex_masks_3_2 : _GEN_35; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_38 = 2'h1 == opidx ? hfutex_masks_1_3 : hfutex_masks_0_3; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_39 = 2'h2 == opidx ? hfutex_masks_2_3 : _GEN_38; // @[NulCtrlMP.scala 166:{48,48}]
  wire [47:0] _GEN_40 = 2'h3 == opidx ? hfutex_masks_3_3 : _GEN_39; // @[NulCtrlMP.scala 166:{48,48}]
  wire  hfutex_hit = _GEN_28 == hfutex_match_reg | _GEN_32 == hfutex_match_reg | _GEN_36 == hfutex_match_reg | _GEN_40
     == hfutex_match_reg; // @[NulCtrlMP.scala 166:79]
  wire  hfutex_hit_set = _GEN_28 == hfutex_set_value | _GEN_32 == hfutex_set_value | _GEN_36 == hfutex_set_value |
    _GEN_40 == hfutex_set_value; // @[NulCtrlMP.scala 167:83]
  reg  send_hear; // @[NulCtrlMP.scala 169:28]
  reg [7:0] uart_buffer; // @[NulCtrlMP.scala 170:30]
  reg [3:0] sleep_cnt; // @[NulCtrlMP.scala 172:28]
  wire [3:0] _sleep_cnt_T_1 = sleep_cnt + 4'h1; // @[NulCtrlMP.scala 174:32]
  wire [4:0] _GEN_41 = sleep_cnt == 4'hf ? 5'h2 : _GEN_20; // @[NulCtrlMP.scala 175:34 176:19]
  wire [4:0] _GEN_43 = state == 5'h1f ? _GEN_41 : _GEN_20; // @[NulCtrlMP.scala 173:33]
  wire  _T_29 = state == 5'h2; // @[NulCtrlMP.scala 180:16]
  wire [4:0] rxop = io_rx_bits[4:0]; // @[NulCtrlMP.scala 183:34]
  wire [2:0] rxoff = io_rx_bits[7:5]; // @[NulCtrlMP.scala 184:35]
  wire [2:0] _GEN_44 = rxop == 5'h0 | rxop == 5'h10 | rxop == 5'h15 ? 3'h4 : 3'h7; // @[NulCtrlMP.scala 208:90 209:23 212:23]
  wire [9:0] _GEN_45 = rxop == 5'h0 | rxop == 5'h10 | rxop == 5'h15 ? 10'h1 : trans_bytes; // @[NulCtrlMP.scala 208:90 210:29 141:30]
  wire [5:0] _GEN_46 = rxop == 5'h0 | rxop == 5'h10 | rxop == 5'h15 ? errno : {{1'd0}, rxop}; // @[NulCtrlMP.scala 144:24 208:90 213:23]
  wire [9:0] _GEN_47 = rxop == 5'hb ? 10'h10 : _GEN_45; // @[NulCtrlMP.scala 206:46 207:29]
  wire [2:0] _GEN_48 = rxop == 5'hb ? 3'h3 : _GEN_44; // @[NulCtrlMP.scala 188:19 206:46]
  wire [5:0] _GEN_49 = rxop == 5'hb ? errno : _GEN_46; // @[NulCtrlMP.scala 144:24 206:46]
  wire [9:0] _GEN_50 = rxop == 5'hd ? 10'hf : _GEN_47; // @[NulCtrlMP.scala 204:45 205:29]
  wire [2:0] _GEN_51 = rxop == 5'hd ? 3'h3 : _GEN_48; // @[NulCtrlMP.scala 188:19 204:45]
  wire [5:0] _GEN_52 = rxop == 5'hd ? errno : _GEN_49; // @[NulCtrlMP.scala 144:24 204:45]
  wire [9:0] _GEN_53 = rxop == 5'h9 | rxop == 5'hf ? 10'hc : _GEN_50; // @[NulCtrlMP.scala 202:69 203:29]
  wire [2:0] _GEN_54 = rxop == 5'h9 | rxop == 5'hf ? 3'h3 : _GEN_51; // @[NulCtrlMP.scala 188:19 202:69]
  wire [5:0] _GEN_55 = rxop == 5'h9 | rxop == 5'hf ? errno : _GEN_52; // @[NulCtrlMP.scala 144:24 202:69]
  wire [9:0] _GEN_56 = rxop == 5'h3 | rxop == 5'h6 ? 10'h9 : _GEN_53; // @[NulCtrlMP.scala 200:68 201:29]
  wire [2:0] _GEN_57 = rxop == 5'h3 | rxop == 5'h6 ? 3'h3 : _GEN_54; // @[NulCtrlMP.scala 188:19 200:68]
  wire [5:0] _GEN_58 = rxop == 5'h3 | rxop == 5'h6 ? errno : _GEN_55; // @[NulCtrlMP.scala 144:24 200:68]
  wire [9:0] _GEN_59 = rxop == 5'h4 | rxop == 5'ha | rxop == 5'h12 ? 10'h8 : _GEN_56; // @[NulCtrlMP.scala 198:94 199:29]
  wire [2:0] _GEN_60 = rxop == 5'h4 | rxop == 5'ha | rxop == 5'h12 ? 3'h3 : _GEN_57; // @[NulCtrlMP.scala 188:19 198:94]
  wire [5:0] _GEN_61 = rxop == 5'h4 | rxop == 5'ha | rxop == 5'h12 ? errno : _GEN_58; // @[NulCtrlMP.scala 144:24 198:94]
  wire [9:0] _GEN_62 = rxop == 5'hc | rxop == 5'he | rxop == 5'h14 ? 10'h7 : _GEN_59; // @[NulCtrlMP.scala 196:93 197:29]
  wire [2:0] _GEN_63 = rxop == 5'hc | rxop == 5'he | rxop == 5'h14 ? 3'h3 : _GEN_60; // @[NulCtrlMP.scala 188:19 196:93]
  wire [5:0] _GEN_64 = rxop == 5'hc | rxop == 5'he | rxop == 5'h14 ? errno : _GEN_61; // @[NulCtrlMP.scala 144:24 196:93]
  wire [9:0] _GEN_65 = rxop == 5'h1e ? 10'h6 : _GEN_62; // @[NulCtrlMP.scala 194:45 195:29]
  wire [2:0] _GEN_66 = rxop == 5'h1e ? 3'h3 : _GEN_63; // @[NulCtrlMP.scala 188:19 194:45]
  wire [5:0] _GEN_67 = rxop == 5'h1e ? errno : _GEN_64; // @[NulCtrlMP.scala 144:24 194:45]
  wire [9:0] _GEN_68 = rxop == 5'h8 ? 10'h4 : _GEN_65; // @[NulCtrlMP.scala 192:46 193:29]
  wire [2:0] _GEN_69 = rxop == 5'h8 ? 3'h3 : _GEN_66; // @[NulCtrlMP.scala 188:19 192:46]
  wire [5:0] _GEN_70 = rxop == 5'h8 ? errno : _GEN_67; // @[NulCtrlMP.scala 144:24 192:46]
  wire [9:0] _GEN_71 = rxop == 5'h1 | rxop == 5'h2 | rxop == 5'h5 | rxop == 5'h7 | rxop == 5'h11 | rxop == 5'h13 ? 10'h2
     : _GEN_68; // @[NulCtrlMP.scala 190:155 191:29]
  wire [2:0] _GEN_72 = rxop == 5'h1 | rxop == 5'h2 | rxop == 5'h5 | rxop == 5'h7 | rxop == 5'h11 | rxop == 5'h13 ? 3'h3
     : _GEN_69; // @[NulCtrlMP.scala 190:155 188:19]
  wire [9:0] _GEN_76 = io_rx_valid ? 10'h1 : trans_pos; // @[NulCtrlMP.scala 182:27 187:23 142:28]
  wire [4:0] _GEN_77 = io_rx_valid ? {{2'd0}, _GEN_72} : _GEN_43; // @[NulCtrlMP.scala 182:27]
  wire [9:0] _GEN_78 = io_rx_valid ? _GEN_71 : trans_bytes; // @[NulCtrlMP.scala 182:27 141:30]
  wire [9:0] _GEN_83 = state == 5'h2 ? _GEN_76 : trans_pos; // @[NulCtrlMP.scala 142:28 180:37]
  wire [4:0] _GEN_84 = state == 5'h2 ? _GEN_77 : _GEN_43; // @[NulCtrlMP.scala 180:37]
  wire [9:0] _GEN_85 = state == 5'h2 ? _GEN_78 : trans_bytes; // @[NulCtrlMP.scala 141:30 180:37]
  wire  _T_66 = state == 5'h3; // @[NulCtrlMP.scala 218:16]
  wire [7:0] _GEN_88 = 4'h1 == trans_pos[3:0] ? io_rx_bits : oparg_1; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_89 = 4'h2 == trans_pos[3:0] ? io_rx_bits : oparg_2; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_90 = 4'h3 == trans_pos[3:0] ? io_rx_bits : oparg_3; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_91 = 4'h4 == trans_pos[3:0] ? io_rx_bits : oparg_4; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_92 = 4'h5 == trans_pos[3:0] ? io_rx_bits : oparg_5; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_93 = 4'h6 == trans_pos[3:0] ? io_rx_bits : oparg_6; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_94 = 4'h7 == trans_pos[3:0] ? io_rx_bits : oparg_7; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_95 = 4'h8 == trans_pos[3:0] ? io_rx_bits : oparg_8; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_96 = 4'h9 == trans_pos[3:0] ? io_rx_bits : oparg_9; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_97 = 4'ha == trans_pos[3:0] ? io_rx_bits : oparg_10; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_98 = 4'hb == trans_pos[3:0] ? io_rx_bits : oparg_11; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_99 = 4'hc == trans_pos[3:0] ? io_rx_bits : oparg_12; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_100 = 4'hd == trans_pos[3:0] ? io_rx_bits : oparg_13; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_101 = 4'he == trans_pos[3:0] ? io_rx_bits : oparg_14; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [7:0] _GEN_102 = 4'hf == trans_pos[3:0] ? io_rx_bits : oparg_15; // @[NulCtrlMP.scala 151:24 221:{30,30}]
  wire [9:0] _T_69 = trans_pos + 10'h1; // @[NulCtrlMP.scala 222:28]
  wire  _T_70 = _T_69 == trans_bytes; // @[NulCtrlMP.scala 222:34]
  wire [9:0] _GEN_103 = _T_69 == trans_bytes ? 10'h0 : _T_69; // @[NulCtrlMP.scala 222:51 223:27 227:27]
  wire [9:0] _GEN_104 = _T_69 == trans_bytes ? 10'h0 : _GEN_85; // @[NulCtrlMP.scala 222:51 224:29]
  wire [4:0] _GEN_105 = _T_69 == trans_bytes ? 5'h4 : _GEN_84; // @[NulCtrlMP.scala 222:51 225:23]
  wire [7:0] _GEN_107 = io_rx_valid ? _GEN_88 : oparg_1; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_108 = io_rx_valid ? _GEN_89 : oparg_2; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_109 = io_rx_valid ? _GEN_90 : oparg_3; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_110 = io_rx_valid ? _GEN_91 : oparg_4; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_111 = io_rx_valid ? _GEN_92 : oparg_5; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_112 = io_rx_valid ? _GEN_93 : oparg_6; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_113 = io_rx_valid ? _GEN_94 : oparg_7; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_114 = io_rx_valid ? _GEN_95 : oparg_8; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_115 = io_rx_valid ? _GEN_96 : oparg_9; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_116 = io_rx_valid ? _GEN_97 : oparg_10; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_117 = io_rx_valid ? _GEN_98 : oparg_11; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_118 = io_rx_valid ? _GEN_99 : oparg_12; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_119 = io_rx_valid ? _GEN_100 : oparg_13; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_120 = io_rx_valid ? _GEN_101 : oparg_14; // @[NulCtrlMP.scala 151:24 220:27]
  wire [7:0] _GEN_121 = io_rx_valid ? _GEN_102 : oparg_15; // @[NulCtrlMP.scala 151:24 220:27]
  wire [9:0] _GEN_122 = io_rx_valid ? _GEN_103 : _GEN_83; // @[NulCtrlMP.scala 220:27]
  wire [9:0] _GEN_123 = io_rx_valid ? _GEN_104 : _GEN_85; // @[NulCtrlMP.scala 220:27]
  wire [4:0] _GEN_124 = io_rx_valid ? _GEN_105 : _GEN_84; // @[NulCtrlMP.scala 220:27]
  wire  _GEN_125 = state == 5'h3 | _T_29; // @[NulCtrlMP.scala 218:36 219:21]
  wire [7:0] _GEN_127 = state == 5'h3 ? _GEN_107 : oparg_1; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_128 = state == 5'h3 ? _GEN_108 : oparg_2; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_129 = state == 5'h3 ? _GEN_109 : oparg_3; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_130 = state == 5'h3 ? _GEN_110 : oparg_4; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_131 = state == 5'h3 ? _GEN_111 : oparg_5; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_132 = state == 5'h3 ? _GEN_112 : oparg_6; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_133 = state == 5'h3 ? _GEN_113 : oparg_7; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_134 = state == 5'h3 ? _GEN_114 : oparg_8; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_135 = state == 5'h3 ? _GEN_115 : oparg_9; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_136 = state == 5'h3 ? _GEN_116 : oparg_10; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_137 = state == 5'h3 ? _GEN_117 : oparg_11; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_138 = state == 5'h3 ? _GEN_118 : oparg_12; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_139 = state == 5'h3 ? _GEN_119 : oparg_13; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_140 = state == 5'h3 ? _GEN_120 : oparg_14; // @[NulCtrlMP.scala 151:24 218:36]
  wire [7:0] _GEN_141 = state == 5'h3 ? _GEN_121 : oparg_15; // @[NulCtrlMP.scala 151:24 218:36]
  wire [9:0] _GEN_142 = state == 5'h3 ? _GEN_122 : _GEN_83; // @[NulCtrlMP.scala 218:36]
  wire [9:0] _GEN_143 = state == 5'h3 ? _GEN_123 : _GEN_85; // @[NulCtrlMP.scala 218:36]
  wire [4:0] _GEN_144 = state == 5'h3 ? _GEN_124 : _GEN_84; // @[NulCtrlMP.scala 218:36]
  wire  _GEN_145 = 2'h0 == opidx; // @[NulCtrlMP.scala 239:{33,33} 44:27]
  wire  _GEN_146 = 2'h1 == opidx; // @[NulCtrlMP.scala 239:{33,33} 44:27]
  wire  _GEN_147 = 2'h2 == opidx; // @[NulCtrlMP.scala 239:{33,33} 44:27]
  wire  _GEN_148 = 2'h3 == opidx; // @[NulCtrlMP.scala 239:{33,33} 44:27]
  wire [1:0] _GEN_149 = 2'h0 == opidx ? 2'h1 : _GEN_21; // @[NulCtrlMP.scala 240:{34,34}]
  wire [1:0] _GEN_150 = 2'h1 == opidx ? 2'h1 : _GEN_22; // @[NulCtrlMP.scala 240:{34,34}]
  wire [1:0] _GEN_151 = 2'h2 == opidx ? 2'h1 : _GEN_23; // @[NulCtrlMP.scala 240:{34,34}]
  wire [1:0] _GEN_152 = 2'h3 == opidx ? 2'h1 : _GEN_24; // @[NulCtrlMP.scala 240:{34,34}]
  wire [1:0] _GEN_158 = 2'h1 == opidx ? cpu_state_1 : cpu_state_0; // @[NulCtrlMP.scala 247:{39,39}]
  wire [1:0] _GEN_159 = 2'h2 == opidx ? cpu_state_2 : _GEN_158; // @[NulCtrlMP.scala 247:{39,39}]
  wire [1:0] _GEN_160 = 2'h3 == opidx ? cpu_state_3 : _GEN_159; // @[NulCtrlMP.scala 247:{39,39}]
  wire [3:0] _GEN_161 = _GEN_160 == 2'h1 | _GEN_160 == 2'h2 ? 4'hb : 4'h5; // @[NulCtrlMP.scala 235:15 247:85 248:27]
  wire [63:0] _GEN_163 = 2'h1 == opidx ? user_clk_1 : user_clk_0; // @[NulCtrlMP.scala 275:{49,49}]
  wire [63:0] _GEN_164 = 2'h2 == opidx ? user_clk_2 : _GEN_163; // @[NulCtrlMP.scala 275:{49,49}]
  wire [63:0] _GEN_165 = 2'h3 == opidx ? user_clk_3 : _GEN_164; // @[NulCtrlMP.scala 275:{49,49}]
  wire [1:0] _GEN_167 = 2'h1 == opidx ? hfutex_pos_1 : hfutex_pos_0; // @[NulCtrlMP.scala 280:{60,60}]
  wire [1:0] _GEN_168 = 2'h2 == opidx ? hfutex_pos_2 : _GEN_167; // @[NulCtrlMP.scala 280:{60,60}]
  wire [1:0] _GEN_169 = 2'h3 == opidx ? hfutex_pos_3 : _GEN_168; // @[NulCtrlMP.scala 280:{60,60}]
  wire [47:0] _GEN_170 = _GEN_145 & 2'h0 == _GEN_169 ? hfutex_set_value : hfutex_masks_0_0; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_171 = _GEN_145 & 2'h1 == _GEN_169 ? hfutex_set_value : hfutex_masks_0_1; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_172 = _GEN_145 & 2'h2 == _GEN_169 ? hfutex_set_value : hfutex_masks_0_2; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_173 = _GEN_145 & 2'h3 == _GEN_169 ? hfutex_set_value : hfutex_masks_0_3; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_174 = _GEN_146 & 2'h0 == _GEN_169 ? hfutex_set_value : hfutex_masks_1_0; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_175 = _GEN_146 & 2'h1 == _GEN_169 ? hfutex_set_value : hfutex_masks_1_1; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_176 = _GEN_146 & 2'h2 == _GEN_169 ? hfutex_set_value : hfutex_masks_1_2; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_177 = _GEN_146 & 2'h3 == _GEN_169 ? hfutex_set_value : hfutex_masks_1_3; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_178 = _GEN_147 & 2'h0 == _GEN_169 ? hfutex_set_value : hfutex_masks_2_0; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_179 = _GEN_147 & 2'h1 == _GEN_169 ? hfutex_set_value : hfutex_masks_2_1; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_180 = _GEN_147 & 2'h2 == _GEN_169 ? hfutex_set_value : hfutex_masks_2_2; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_181 = _GEN_147 & 2'h3 == _GEN_169 ? hfutex_set_value : hfutex_masks_2_3; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_182 = _GEN_148 & 2'h0 == _GEN_169 ? hfutex_set_value : hfutex_masks_3_0; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_183 = _GEN_148 & 2'h1 == _GEN_169 ? hfutex_set_value : hfutex_masks_3_1; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_184 = _GEN_148 & 2'h2 == _GEN_169 ? hfutex_set_value : hfutex_masks_3_2; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [47:0] _GEN_185 = _GEN_148 & 2'h3 == _GEN_169 ? hfutex_set_value : hfutex_masks_3_3; // @[NulCtrlMP.scala 162:31 280:{60,60}]
  wire [1:0] _hfutex_pos_T_2 = _GEN_169 + 2'h1; // @[NulCtrlMP.scala 281:96]
  wire [1:0] _hfutex_pos_T_3 = _GEN_169 == 2'h3 ? 2'h0 : _hfutex_pos_T_2; // @[NulCtrlMP.scala 281:45]
  wire [1:0] _GEN_186 = 2'h0 == opidx ? _hfutex_pos_T_3 : hfutex_pos_0; // @[NulCtrlMP.scala 163:29 281:{39,39}]
  wire [1:0] _GEN_187 = 2'h1 == opidx ? _hfutex_pos_T_3 : hfutex_pos_1; // @[NulCtrlMP.scala 163:29 281:{39,39}]
  wire [1:0] _GEN_188 = 2'h2 == opidx ? _hfutex_pos_T_3 : hfutex_pos_2; // @[NulCtrlMP.scala 163:29 281:{39,39}]
  wire [1:0] _GEN_189 = 2'h3 == opidx ? _hfutex_pos_T_3 : hfutex_pos_3; // @[NulCtrlMP.scala 163:29 281:{39,39}]
  wire [47:0] _GEN_190 = ~hfutex_hit_set ? _GEN_170 : hfutex_masks_0_0; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_191 = ~hfutex_hit_set ? _GEN_171 : hfutex_masks_0_1; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_192 = ~hfutex_hit_set ? _GEN_172 : hfutex_masks_0_2; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_193 = ~hfutex_hit_set ? _GEN_173 : hfutex_masks_0_3; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_194 = ~hfutex_hit_set ? _GEN_174 : hfutex_masks_1_0; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_195 = ~hfutex_hit_set ? _GEN_175 : hfutex_masks_1_1; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_196 = ~hfutex_hit_set ? _GEN_176 : hfutex_masks_1_2; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_197 = ~hfutex_hit_set ? _GEN_177 : hfutex_masks_1_3; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_198 = ~hfutex_hit_set ? _GEN_178 : hfutex_masks_2_0; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_199 = ~hfutex_hit_set ? _GEN_179 : hfutex_masks_2_1; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_200 = ~hfutex_hit_set ? _GEN_180 : hfutex_masks_2_2; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_201 = ~hfutex_hit_set ? _GEN_181 : hfutex_masks_2_3; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_202 = ~hfutex_hit_set ? _GEN_182 : hfutex_masks_3_0; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_203 = ~hfutex_hit_set ? _GEN_183 : hfutex_masks_3_1; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_204 = ~hfutex_hit_set ? _GEN_184 : hfutex_masks_3_2; // @[NulCtrlMP.scala 162:31 279:39]
  wire [47:0] _GEN_205 = ~hfutex_hit_set ? _GEN_185 : hfutex_masks_3_3; // @[NulCtrlMP.scala 162:31 279:39]
  wire [1:0] _GEN_206 = ~hfutex_hit_set ? _GEN_186 : hfutex_pos_0; // @[NulCtrlMP.scala 163:29 279:39]
  wire [1:0] _GEN_207 = ~hfutex_hit_set ? _GEN_187 : hfutex_pos_1; // @[NulCtrlMP.scala 163:29 279:39]
  wire [1:0] _GEN_208 = ~hfutex_hit_set ? _GEN_188 : hfutex_pos_2; // @[NulCtrlMP.scala 163:29 279:39]
  wire [1:0] _GEN_209 = ~hfutex_hit_set ? _GEN_189 : hfutex_pos_3; // @[NulCtrlMP.scala 163:29 279:39]
  wire [47:0] _GEN_210 = 2'h0 == opidx ? 48'h0 : hfutex_masks_0_0; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_211 = 2'h1 == opidx ? 48'h0 : hfutex_masks_1_0; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_212 = 2'h2 == opidx ? 48'h0 : hfutex_masks_2_0; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_213 = 2'h3 == opidx ? 48'h0 : hfutex_masks_3_0; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_214 = 2'h0 == opidx ? 48'h0 : hfutex_masks_0_1; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_215 = 2'h1 == opidx ? 48'h0 : hfutex_masks_1_1; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_216 = 2'h2 == opidx ? 48'h0 : hfutex_masks_2_1; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_217 = 2'h3 == opidx ? 48'h0 : hfutex_masks_3_1; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_218 = 2'h0 == opidx ? 48'h0 : hfutex_masks_0_2; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_219 = 2'h1 == opidx ? 48'h0 : hfutex_masks_1_2; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_220 = 2'h2 == opidx ? 48'h0 : hfutex_masks_2_2; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_221 = 2'h3 == opidx ? 48'h0 : hfutex_masks_3_2; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_222 = 2'h0 == opidx ? 48'h0 : hfutex_masks_0_3; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_223 = 2'h1 == opidx ? 48'h0 : hfutex_masks_1_3; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_224 = 2'h2 == opidx ? 48'h0 : hfutex_masks_2_3; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [47:0] _GEN_225 = 2'h3 == opidx ? 48'h0 : hfutex_masks_3_3; // @[NulCtrlMP.scala 162:31 286:{44,44}]
  wire [4:0] _GEN_226 = 5'h15 == opcode ? 5'h19 : 5'h5; // @[NulCtrlMP.scala 235:15 236:24 291:21]
  wire  _GEN_227 = 5'h15 == opcode ? 1'h0 : send_hear; // @[NulCtrlMP.scala 236:24 292:25 169:28]
  wire [4:0] _GEN_228 = 5'h1e == opcode ? 5'h17 : _GEN_226; // @[NulCtrlMP.scala 236:24 289:36]
  wire  _GEN_229 = 5'h1e == opcode ? send_hear : _GEN_227; // @[NulCtrlMP.scala 236:24 169:28]
  wire [47:0] _GEN_230 = 5'h13 == opcode ? _GEN_210 : hfutex_masks_0_0; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_231 = 5'h13 == opcode ? _GEN_211 : hfutex_masks_1_0; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_232 = 5'h13 == opcode ? _GEN_212 : hfutex_masks_2_0; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_233 = 5'h13 == opcode ? _GEN_213 : hfutex_masks_3_0; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_234 = 5'h13 == opcode ? _GEN_214 : hfutex_masks_0_1; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_235 = 5'h13 == opcode ? _GEN_215 : hfutex_masks_1_1; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_236 = 5'h13 == opcode ? _GEN_216 : hfutex_masks_2_1; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_237 = 5'h13 == opcode ? _GEN_217 : hfutex_masks_3_1; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_238 = 5'h13 == opcode ? _GEN_218 : hfutex_masks_0_2; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_239 = 5'h13 == opcode ? _GEN_219 : hfutex_masks_1_2; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_240 = 5'h13 == opcode ? _GEN_220 : hfutex_masks_2_2; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_241 = 5'h13 == opcode ? _GEN_221 : hfutex_masks_3_2; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_242 = 5'h13 == opcode ? _GEN_222 : hfutex_masks_0_3; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_243 = 5'h13 == opcode ? _GEN_223 : hfutex_masks_1_3; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_244 = 5'h13 == opcode ? _GEN_224 : hfutex_masks_2_3; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_245 = 5'h13 == opcode ? _GEN_225 : hfutex_masks_3_3; // @[NulCtrlMP.scala 236:24 162:31]
  wire [4:0] _GEN_246 = 5'h13 == opcode ? 5'h5 : _GEN_228; // @[NulCtrlMP.scala 235:15 236:24]
  wire  _GEN_247 = 5'h13 == opcode ? send_hear : _GEN_229; // @[NulCtrlMP.scala 236:24 169:28]
  wire [47:0] _GEN_248 = 5'h12 == opcode ? _GEN_190 : _GEN_230; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_249 = 5'h12 == opcode ? _GEN_191 : _GEN_234; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_250 = 5'h12 == opcode ? _GEN_192 : _GEN_238; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_251 = 5'h12 == opcode ? _GEN_193 : _GEN_242; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_252 = 5'h12 == opcode ? _GEN_194 : _GEN_231; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_253 = 5'h12 == opcode ? _GEN_195 : _GEN_235; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_254 = 5'h12 == opcode ? _GEN_196 : _GEN_239; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_255 = 5'h12 == opcode ? _GEN_197 : _GEN_243; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_256 = 5'h12 == opcode ? _GEN_198 : _GEN_232; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_257 = 5'h12 == opcode ? _GEN_199 : _GEN_236; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_258 = 5'h12 == opcode ? _GEN_200 : _GEN_240; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_259 = 5'h12 == opcode ? _GEN_201 : _GEN_244; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_260 = 5'h12 == opcode ? _GEN_202 : _GEN_233; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_261 = 5'h12 == opcode ? _GEN_203 : _GEN_237; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_262 = 5'h12 == opcode ? _GEN_204 : _GEN_241; // @[NulCtrlMP.scala 236:24]
  wire [47:0] _GEN_263 = 5'h12 == opcode ? _GEN_205 : _GEN_245; // @[NulCtrlMP.scala 236:24]
  wire [1:0] _GEN_264 = 5'h12 == opcode ? _GEN_206 : hfutex_pos_0; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_265 = 5'h12 == opcode ? _GEN_207 : hfutex_pos_1; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_266 = 5'h12 == opcode ? _GEN_208 : hfutex_pos_2; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_267 = 5'h12 == opcode ? _GEN_209 : hfutex_pos_3; // @[NulCtrlMP.scala 236:24 163:29]
  wire [4:0] _GEN_268 = 5'h12 == opcode ? 5'h5 : _GEN_246; // @[NulCtrlMP.scala 235:15 236:24]
  wire  _GEN_269 = 5'h12 == opcode ? send_hear : _GEN_247; // @[NulCtrlMP.scala 236:24 169:28]
  wire [7:0] _GEN_270 = 5'h11 == opcode ? _GEN_165[7:0] : retarg_0; // @[NulCtrlMP.scala 236:24 152:25 275:31]
  wire [7:0] _GEN_271 = 5'h11 == opcode ? _GEN_165[15:8] : retarg_1; // @[NulCtrlMP.scala 236:24 152:25 275:31]
  wire [7:0] _GEN_272 = 5'h11 == opcode ? _GEN_165[23:16] : retarg_2; // @[NulCtrlMP.scala 236:24 152:25 275:31]
  wire [7:0] _GEN_273 = 5'h11 == opcode ? _GEN_165[31:24] : retarg_3; // @[NulCtrlMP.scala 236:24 152:25 275:31]
  wire [7:0] _GEN_274 = 5'h11 == opcode ? _GEN_165[39:32] : retarg_4; // @[NulCtrlMP.scala 236:24 152:25 275:31]
  wire [7:0] _GEN_275 = 5'h11 == opcode ? _GEN_165[47:40] : retarg_5; // @[NulCtrlMP.scala 236:24 152:25 275:31]
  wire [7:0] _GEN_276 = 5'h11 == opcode ? _GEN_165[55:48] : retarg_6; // @[NulCtrlMP.scala 236:24 152:25 275:31]
  wire [7:0] _GEN_277 = 5'h11 == opcode ? _GEN_165[63:56] : retarg_7; // @[NulCtrlMP.scala 236:24 152:25 275:31]
  wire [47:0] _GEN_278 = 5'h11 == opcode ? hfutex_masks_0_0 : _GEN_248; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_279 = 5'h11 == opcode ? hfutex_masks_0_1 : _GEN_249; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_280 = 5'h11 == opcode ? hfutex_masks_0_2 : _GEN_250; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_281 = 5'h11 == opcode ? hfutex_masks_0_3 : _GEN_251; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_282 = 5'h11 == opcode ? hfutex_masks_1_0 : _GEN_252; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_283 = 5'h11 == opcode ? hfutex_masks_1_1 : _GEN_253; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_284 = 5'h11 == opcode ? hfutex_masks_1_2 : _GEN_254; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_285 = 5'h11 == opcode ? hfutex_masks_1_3 : _GEN_255; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_286 = 5'h11 == opcode ? hfutex_masks_2_0 : _GEN_256; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_287 = 5'h11 == opcode ? hfutex_masks_2_1 : _GEN_257; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_288 = 5'h11 == opcode ? hfutex_masks_2_2 : _GEN_258; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_289 = 5'h11 == opcode ? hfutex_masks_2_3 : _GEN_259; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_290 = 5'h11 == opcode ? hfutex_masks_3_0 : _GEN_260; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_291 = 5'h11 == opcode ? hfutex_masks_3_1 : _GEN_261; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_292 = 5'h11 == opcode ? hfutex_masks_3_2 : _GEN_262; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_293 = 5'h11 == opcode ? hfutex_masks_3_3 : _GEN_263; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_294 = 5'h11 == opcode ? hfutex_pos_0 : _GEN_264; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_295 = 5'h11 == opcode ? hfutex_pos_1 : _GEN_265; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_296 = 5'h11 == opcode ? hfutex_pos_2 : _GEN_266; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_297 = 5'h11 == opcode ? hfutex_pos_3 : _GEN_267; // @[NulCtrlMP.scala 236:24 163:29]
  wire [4:0] _GEN_298 = 5'h11 == opcode ? 5'h5 : _GEN_268; // @[NulCtrlMP.scala 235:15 236:24]
  wire  _GEN_299 = 5'h11 == opcode ? send_hear : _GEN_269; // @[NulCtrlMP.scala 236:24 169:28]
  wire [7:0] _GEN_300 = 5'h10 == opcode ? global_clk[7:0] : _GEN_270; // @[NulCtrlMP.scala 236:24 270:31]
  wire [7:0] _GEN_301 = 5'h10 == opcode ? global_clk[15:8] : _GEN_271; // @[NulCtrlMP.scala 236:24 270:31]
  wire [7:0] _GEN_302 = 5'h10 == opcode ? global_clk[23:16] : _GEN_272; // @[NulCtrlMP.scala 236:24 270:31]
  wire [7:0] _GEN_303 = 5'h10 == opcode ? global_clk[31:24] : _GEN_273; // @[NulCtrlMP.scala 236:24 270:31]
  wire [7:0] _GEN_304 = 5'h10 == opcode ? global_clk[39:32] : _GEN_274; // @[NulCtrlMP.scala 236:24 270:31]
  wire [7:0] _GEN_305 = 5'h10 == opcode ? global_clk[47:40] : _GEN_275; // @[NulCtrlMP.scala 236:24 270:31]
  wire [7:0] _GEN_306 = 5'h10 == opcode ? global_clk[55:48] : _GEN_276; // @[NulCtrlMP.scala 236:24 270:31]
  wire [7:0] _GEN_307 = 5'h10 == opcode ? global_clk[63:56] : _GEN_277; // @[NulCtrlMP.scala 236:24 270:31]
  wire [47:0] _GEN_308 = 5'h10 == opcode ? hfutex_masks_0_0 : _GEN_278; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_309 = 5'h10 == opcode ? hfutex_masks_0_1 : _GEN_279; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_310 = 5'h10 == opcode ? hfutex_masks_0_2 : _GEN_280; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_311 = 5'h10 == opcode ? hfutex_masks_0_3 : _GEN_281; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_312 = 5'h10 == opcode ? hfutex_masks_1_0 : _GEN_282; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_313 = 5'h10 == opcode ? hfutex_masks_1_1 : _GEN_283; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_314 = 5'h10 == opcode ? hfutex_masks_1_2 : _GEN_284; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_315 = 5'h10 == opcode ? hfutex_masks_1_3 : _GEN_285; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_316 = 5'h10 == opcode ? hfutex_masks_2_0 : _GEN_286; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_317 = 5'h10 == opcode ? hfutex_masks_2_1 : _GEN_287; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_318 = 5'h10 == opcode ? hfutex_masks_2_2 : _GEN_288; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_319 = 5'h10 == opcode ? hfutex_masks_2_3 : _GEN_289; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_320 = 5'h10 == opcode ? hfutex_masks_3_0 : _GEN_290; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_321 = 5'h10 == opcode ? hfutex_masks_3_1 : _GEN_291; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_322 = 5'h10 == opcode ? hfutex_masks_3_2 : _GEN_292; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_323 = 5'h10 == opcode ? hfutex_masks_3_3 : _GEN_293; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_324 = 5'h10 == opcode ? hfutex_pos_0 : _GEN_294; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_325 = 5'h10 == opcode ? hfutex_pos_1 : _GEN_295; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_326 = 5'h10 == opcode ? hfutex_pos_2 : _GEN_296; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_327 = 5'h10 == opcode ? hfutex_pos_3 : _GEN_297; // @[NulCtrlMP.scala 236:24 163:29]
  wire [4:0] _GEN_328 = 5'h10 == opcode ? 5'h5 : _GEN_298; // @[NulCtrlMP.scala 235:15 236:24]
  wire  _GEN_329 = 5'h10 == opcode ? send_hear : _GEN_299; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_330 = 5'hf == opcode ? 5'h15 : _GEN_328; // @[NulCtrlMP.scala 236:24 267:36]
  wire [7:0] _GEN_331 = 5'hf == opcode ? retarg_0 : _GEN_300; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_332 = 5'hf == opcode ? retarg_1 : _GEN_301; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_333 = 5'hf == opcode ? retarg_2 : _GEN_302; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_334 = 5'hf == opcode ? retarg_3 : _GEN_303; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_335 = 5'hf == opcode ? retarg_4 : _GEN_304; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_336 = 5'hf == opcode ? retarg_5 : _GEN_305; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_337 = 5'hf == opcode ? retarg_6 : _GEN_306; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_338 = 5'hf == opcode ? retarg_7 : _GEN_307; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_339 = 5'hf == opcode ? hfutex_masks_0_0 : _GEN_308; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_340 = 5'hf == opcode ? hfutex_masks_0_1 : _GEN_309; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_341 = 5'hf == opcode ? hfutex_masks_0_2 : _GEN_310; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_342 = 5'hf == opcode ? hfutex_masks_0_3 : _GEN_311; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_343 = 5'hf == opcode ? hfutex_masks_1_0 : _GEN_312; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_344 = 5'hf == opcode ? hfutex_masks_1_1 : _GEN_313; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_345 = 5'hf == opcode ? hfutex_masks_1_2 : _GEN_314; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_346 = 5'hf == opcode ? hfutex_masks_1_3 : _GEN_315; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_347 = 5'hf == opcode ? hfutex_masks_2_0 : _GEN_316; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_348 = 5'hf == opcode ? hfutex_masks_2_1 : _GEN_317; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_349 = 5'hf == opcode ? hfutex_masks_2_2 : _GEN_318; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_350 = 5'hf == opcode ? hfutex_masks_2_3 : _GEN_319; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_351 = 5'hf == opcode ? hfutex_masks_3_0 : _GEN_320; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_352 = 5'hf == opcode ? hfutex_masks_3_1 : _GEN_321; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_353 = 5'hf == opcode ? hfutex_masks_3_2 : _GEN_322; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_354 = 5'hf == opcode ? hfutex_masks_3_3 : _GEN_323; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_355 = 5'hf == opcode ? hfutex_pos_0 : _GEN_324; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_356 = 5'hf == opcode ? hfutex_pos_1 : _GEN_325; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_357 = 5'hf == opcode ? hfutex_pos_2 : _GEN_326; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_358 = 5'hf == opcode ? hfutex_pos_3 : _GEN_327; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_359 = 5'hf == opcode ? send_hear : _GEN_329; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_360 = 5'he == opcode ? 5'h14 : _GEN_330; // @[NulCtrlMP.scala 236:24 266:36]
  wire [7:0] _GEN_361 = 5'he == opcode ? retarg_0 : _GEN_331; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_362 = 5'he == opcode ? retarg_1 : _GEN_332; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_363 = 5'he == opcode ? retarg_2 : _GEN_333; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_364 = 5'he == opcode ? retarg_3 : _GEN_334; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_365 = 5'he == opcode ? retarg_4 : _GEN_335; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_366 = 5'he == opcode ? retarg_5 : _GEN_336; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_367 = 5'he == opcode ? retarg_6 : _GEN_337; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_368 = 5'he == opcode ? retarg_7 : _GEN_338; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_369 = 5'he == opcode ? hfutex_masks_0_0 : _GEN_339; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_370 = 5'he == opcode ? hfutex_masks_0_1 : _GEN_340; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_371 = 5'he == opcode ? hfutex_masks_0_2 : _GEN_341; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_372 = 5'he == opcode ? hfutex_masks_0_3 : _GEN_342; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_373 = 5'he == opcode ? hfutex_masks_1_0 : _GEN_343; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_374 = 5'he == opcode ? hfutex_masks_1_1 : _GEN_344; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_375 = 5'he == opcode ? hfutex_masks_1_2 : _GEN_345; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_376 = 5'he == opcode ? hfutex_masks_1_3 : _GEN_346; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_377 = 5'he == opcode ? hfutex_masks_2_0 : _GEN_347; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_378 = 5'he == opcode ? hfutex_masks_2_1 : _GEN_348; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_379 = 5'he == opcode ? hfutex_masks_2_2 : _GEN_349; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_380 = 5'he == opcode ? hfutex_masks_2_3 : _GEN_350; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_381 = 5'he == opcode ? hfutex_masks_3_0 : _GEN_351; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_382 = 5'he == opcode ? hfutex_masks_3_1 : _GEN_352; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_383 = 5'he == opcode ? hfutex_masks_3_2 : _GEN_353; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_384 = 5'he == opcode ? hfutex_masks_3_3 : _GEN_354; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_385 = 5'he == opcode ? hfutex_pos_0 : _GEN_355; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_386 = 5'he == opcode ? hfutex_pos_1 : _GEN_356; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_387 = 5'he == opcode ? hfutex_pos_2 : _GEN_357; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_388 = 5'he == opcode ? hfutex_pos_3 : _GEN_358; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_389 = 5'he == opcode ? send_hear : _GEN_359; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_390 = 5'h14 == opcode ? 5'h13 : _GEN_360; // @[NulCtrlMP.scala 236:24 261:23]
  wire [7:0] _GEN_391 = 5'h14 == opcode ? 8'h0 : _GEN_133; // @[NulCtrlMP.scala 236:24 263:34]
  wire [7:0] _GEN_392 = 5'h14 == opcode ? 8'h0 : _GEN_134; // @[NulCtrlMP.scala 236:24 263:34]
  wire [7:0] _GEN_393 = 5'h14 == opcode ? 8'h0 : _GEN_135; // @[NulCtrlMP.scala 236:24 263:34]
  wire [7:0] _GEN_394 = 5'h14 == opcode ? 8'h0 : _GEN_136; // @[NulCtrlMP.scala 236:24 263:34]
  wire [7:0] _GEN_395 = 5'h14 == opcode ? 8'h0 : _GEN_137; // @[NulCtrlMP.scala 236:24 263:34]
  wire [7:0] _GEN_396 = 5'h14 == opcode ? 8'h0 : _GEN_138; // @[NulCtrlMP.scala 236:24 263:34]
  wire [7:0] _GEN_397 = 5'h14 == opcode ? 8'h0 : _GEN_139; // @[NulCtrlMP.scala 236:24 263:34]
  wire [7:0] _GEN_398 = 5'h14 == opcode ? 8'h0 : _GEN_140; // @[NulCtrlMP.scala 236:24 263:34]
  wire [7:0] _GEN_399 = 5'h14 == opcode ? retarg_0 : _GEN_361; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_400 = 5'h14 == opcode ? retarg_1 : _GEN_362; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_401 = 5'h14 == opcode ? retarg_2 : _GEN_363; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_402 = 5'h14 == opcode ? retarg_3 : _GEN_364; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_403 = 5'h14 == opcode ? retarg_4 : _GEN_365; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_404 = 5'h14 == opcode ? retarg_5 : _GEN_366; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_405 = 5'h14 == opcode ? retarg_6 : _GEN_367; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_406 = 5'h14 == opcode ? retarg_7 : _GEN_368; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_407 = 5'h14 == opcode ? hfutex_masks_0_0 : _GEN_369; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_408 = 5'h14 == opcode ? hfutex_masks_0_1 : _GEN_370; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_409 = 5'h14 == opcode ? hfutex_masks_0_2 : _GEN_371; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_410 = 5'h14 == opcode ? hfutex_masks_0_3 : _GEN_372; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_411 = 5'h14 == opcode ? hfutex_masks_1_0 : _GEN_373; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_412 = 5'h14 == opcode ? hfutex_masks_1_1 : _GEN_374; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_413 = 5'h14 == opcode ? hfutex_masks_1_2 : _GEN_375; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_414 = 5'h14 == opcode ? hfutex_masks_1_3 : _GEN_376; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_415 = 5'h14 == opcode ? hfutex_masks_2_0 : _GEN_377; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_416 = 5'h14 == opcode ? hfutex_masks_2_1 : _GEN_378; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_417 = 5'h14 == opcode ? hfutex_masks_2_2 : _GEN_379; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_418 = 5'h14 == opcode ? hfutex_masks_2_3 : _GEN_380; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_419 = 5'h14 == opcode ? hfutex_masks_3_0 : _GEN_381; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_420 = 5'h14 == opcode ? hfutex_masks_3_1 : _GEN_382; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_421 = 5'h14 == opcode ? hfutex_masks_3_2 : _GEN_383; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_422 = 5'h14 == opcode ? hfutex_masks_3_3 : _GEN_384; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_423 = 5'h14 == opcode ? hfutex_pos_0 : _GEN_385; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_424 = 5'h14 == opcode ? hfutex_pos_1 : _GEN_386; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_425 = 5'h14 == opcode ? hfutex_pos_2 : _GEN_387; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_426 = 5'h14 == opcode ? hfutex_pos_3 : _GEN_388; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_427 = 5'h14 == opcode ? send_hear : _GEN_389; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_428 = 5'hd == opcode ? 5'h13 : _GEN_390; // @[NulCtrlMP.scala 236:24 259:36]
  wire [7:0] _GEN_429 = 5'hd == opcode ? _GEN_133 : _GEN_391; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_430 = 5'hd == opcode ? _GEN_134 : _GEN_392; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_431 = 5'hd == opcode ? _GEN_135 : _GEN_393; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_432 = 5'hd == opcode ? _GEN_136 : _GEN_394; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_433 = 5'hd == opcode ? _GEN_137 : _GEN_395; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_434 = 5'hd == opcode ? _GEN_138 : _GEN_396; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_435 = 5'hd == opcode ? _GEN_139 : _GEN_397; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_436 = 5'hd == opcode ? _GEN_140 : _GEN_398; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_437 = 5'hd == opcode ? retarg_0 : _GEN_399; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_438 = 5'hd == opcode ? retarg_1 : _GEN_400; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_439 = 5'hd == opcode ? retarg_2 : _GEN_401; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_440 = 5'hd == opcode ? retarg_3 : _GEN_402; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_441 = 5'hd == opcode ? retarg_4 : _GEN_403; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_442 = 5'hd == opcode ? retarg_5 : _GEN_404; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_443 = 5'hd == opcode ? retarg_6 : _GEN_405; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_444 = 5'hd == opcode ? retarg_7 : _GEN_406; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_445 = 5'hd == opcode ? hfutex_masks_0_0 : _GEN_407; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_446 = 5'hd == opcode ? hfutex_masks_0_1 : _GEN_408; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_447 = 5'hd == opcode ? hfutex_masks_0_2 : _GEN_409; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_448 = 5'hd == opcode ? hfutex_masks_0_3 : _GEN_410; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_449 = 5'hd == opcode ? hfutex_masks_1_0 : _GEN_411; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_450 = 5'hd == opcode ? hfutex_masks_1_1 : _GEN_412; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_451 = 5'hd == opcode ? hfutex_masks_1_2 : _GEN_413; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_452 = 5'hd == opcode ? hfutex_masks_1_3 : _GEN_414; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_453 = 5'hd == opcode ? hfutex_masks_2_0 : _GEN_415; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_454 = 5'hd == opcode ? hfutex_masks_2_1 : _GEN_416; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_455 = 5'hd == opcode ? hfutex_masks_2_2 : _GEN_417; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_456 = 5'hd == opcode ? hfutex_masks_2_3 : _GEN_418; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_457 = 5'hd == opcode ? hfutex_masks_3_0 : _GEN_419; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_458 = 5'hd == opcode ? hfutex_masks_3_1 : _GEN_420; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_459 = 5'hd == opcode ? hfutex_masks_3_2 : _GEN_421; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_460 = 5'hd == opcode ? hfutex_masks_3_3 : _GEN_422; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_461 = 5'hd == opcode ? hfutex_pos_0 : _GEN_423; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_462 = 5'hd == opcode ? hfutex_pos_1 : _GEN_424; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_463 = 5'hd == opcode ? hfutex_pos_2 : _GEN_425; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_464 = 5'hd == opcode ? hfutex_pos_3 : _GEN_426; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_465 = 5'hd == opcode ? send_hear : _GEN_427; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_466 = 5'hc == opcode ? 5'h12 : _GEN_428; // @[NulCtrlMP.scala 236:24 258:36]
  wire [7:0] _GEN_467 = 5'hc == opcode ? _GEN_133 : _GEN_429; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_468 = 5'hc == opcode ? _GEN_134 : _GEN_430; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_469 = 5'hc == opcode ? _GEN_135 : _GEN_431; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_470 = 5'hc == opcode ? _GEN_136 : _GEN_432; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_471 = 5'hc == opcode ? _GEN_137 : _GEN_433; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_472 = 5'hc == opcode ? _GEN_138 : _GEN_434; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_473 = 5'hc == opcode ? _GEN_139 : _GEN_435; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_474 = 5'hc == opcode ? _GEN_140 : _GEN_436; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_475 = 5'hc == opcode ? retarg_0 : _GEN_437; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_476 = 5'hc == opcode ? retarg_1 : _GEN_438; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_477 = 5'hc == opcode ? retarg_2 : _GEN_439; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_478 = 5'hc == opcode ? retarg_3 : _GEN_440; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_479 = 5'hc == opcode ? retarg_4 : _GEN_441; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_480 = 5'hc == opcode ? retarg_5 : _GEN_442; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_481 = 5'hc == opcode ? retarg_6 : _GEN_443; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_482 = 5'hc == opcode ? retarg_7 : _GEN_444; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_483 = 5'hc == opcode ? hfutex_masks_0_0 : _GEN_445; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_484 = 5'hc == opcode ? hfutex_masks_0_1 : _GEN_446; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_485 = 5'hc == opcode ? hfutex_masks_0_2 : _GEN_447; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_486 = 5'hc == opcode ? hfutex_masks_0_3 : _GEN_448; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_487 = 5'hc == opcode ? hfutex_masks_1_0 : _GEN_449; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_488 = 5'hc == opcode ? hfutex_masks_1_1 : _GEN_450; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_489 = 5'hc == opcode ? hfutex_masks_1_2 : _GEN_451; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_490 = 5'hc == opcode ? hfutex_masks_1_3 : _GEN_452; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_491 = 5'hc == opcode ? hfutex_masks_2_0 : _GEN_453; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_492 = 5'hc == opcode ? hfutex_masks_2_1 : _GEN_454; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_493 = 5'hc == opcode ? hfutex_masks_2_2 : _GEN_455; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_494 = 5'hc == opcode ? hfutex_masks_2_3 : _GEN_456; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_495 = 5'hc == opcode ? hfutex_masks_3_0 : _GEN_457; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_496 = 5'hc == opcode ? hfutex_masks_3_1 : _GEN_458; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_497 = 5'hc == opcode ? hfutex_masks_3_2 : _GEN_459; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_498 = 5'hc == opcode ? hfutex_masks_3_3 : _GEN_460; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_499 = 5'hc == opcode ? hfutex_pos_0 : _GEN_461; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_500 = 5'hc == opcode ? hfutex_pos_1 : _GEN_462; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_501 = 5'hc == opcode ? hfutex_pos_2 : _GEN_463; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_502 = 5'hc == opcode ? hfutex_pos_3 : _GEN_464; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_503 = 5'hc == opcode ? send_hear : _GEN_465; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_504 = 5'hb == opcode ? 5'h11 : _GEN_466; // @[NulCtrlMP.scala 236:24 257:37]
  wire [7:0] _GEN_505 = 5'hb == opcode ? _GEN_133 : _GEN_467; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_506 = 5'hb == opcode ? _GEN_134 : _GEN_468; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_507 = 5'hb == opcode ? _GEN_135 : _GEN_469; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_508 = 5'hb == opcode ? _GEN_136 : _GEN_470; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_509 = 5'hb == opcode ? _GEN_137 : _GEN_471; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_510 = 5'hb == opcode ? _GEN_138 : _GEN_472; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_511 = 5'hb == opcode ? _GEN_139 : _GEN_473; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_512 = 5'hb == opcode ? _GEN_140 : _GEN_474; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_513 = 5'hb == opcode ? retarg_0 : _GEN_475; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_514 = 5'hb == opcode ? retarg_1 : _GEN_476; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_515 = 5'hb == opcode ? retarg_2 : _GEN_477; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_516 = 5'hb == opcode ? retarg_3 : _GEN_478; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_517 = 5'hb == opcode ? retarg_4 : _GEN_479; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_518 = 5'hb == opcode ? retarg_5 : _GEN_480; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_519 = 5'hb == opcode ? retarg_6 : _GEN_481; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_520 = 5'hb == opcode ? retarg_7 : _GEN_482; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_521 = 5'hb == opcode ? hfutex_masks_0_0 : _GEN_483; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_522 = 5'hb == opcode ? hfutex_masks_0_1 : _GEN_484; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_523 = 5'hb == opcode ? hfutex_masks_0_2 : _GEN_485; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_524 = 5'hb == opcode ? hfutex_masks_0_3 : _GEN_486; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_525 = 5'hb == opcode ? hfutex_masks_1_0 : _GEN_487; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_526 = 5'hb == opcode ? hfutex_masks_1_1 : _GEN_488; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_527 = 5'hb == opcode ? hfutex_masks_1_2 : _GEN_489; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_528 = 5'hb == opcode ? hfutex_masks_1_3 : _GEN_490; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_529 = 5'hb == opcode ? hfutex_masks_2_0 : _GEN_491; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_530 = 5'hb == opcode ? hfutex_masks_2_1 : _GEN_492; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_531 = 5'hb == opcode ? hfutex_masks_2_2 : _GEN_493; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_532 = 5'hb == opcode ? hfutex_masks_2_3 : _GEN_494; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_533 = 5'hb == opcode ? hfutex_masks_3_0 : _GEN_495; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_534 = 5'hb == opcode ? hfutex_masks_3_1 : _GEN_496; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_535 = 5'hb == opcode ? hfutex_masks_3_2 : _GEN_497; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_536 = 5'hb == opcode ? hfutex_masks_3_3 : _GEN_498; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_537 = 5'hb == opcode ? hfutex_pos_0 : _GEN_499; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_538 = 5'hb == opcode ? hfutex_pos_1 : _GEN_500; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_539 = 5'hb == opcode ? hfutex_pos_2 : _GEN_501; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_540 = 5'hb == opcode ? hfutex_pos_3 : _GEN_502; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_541 = 5'hb == opcode ? send_hear : _GEN_503; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_542 = 5'ha == opcode ? 5'h10 : _GEN_504; // @[NulCtrlMP.scala 236:24 256:37]
  wire [7:0] _GEN_543 = 5'ha == opcode ? _GEN_133 : _GEN_505; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_544 = 5'ha == opcode ? _GEN_134 : _GEN_506; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_545 = 5'ha == opcode ? _GEN_135 : _GEN_507; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_546 = 5'ha == opcode ? _GEN_136 : _GEN_508; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_547 = 5'ha == opcode ? _GEN_137 : _GEN_509; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_548 = 5'ha == opcode ? _GEN_138 : _GEN_510; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_549 = 5'ha == opcode ? _GEN_139 : _GEN_511; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_550 = 5'ha == opcode ? _GEN_140 : _GEN_512; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_551 = 5'ha == opcode ? retarg_0 : _GEN_513; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_552 = 5'ha == opcode ? retarg_1 : _GEN_514; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_553 = 5'ha == opcode ? retarg_2 : _GEN_515; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_554 = 5'ha == opcode ? retarg_3 : _GEN_516; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_555 = 5'ha == opcode ? retarg_4 : _GEN_517; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_556 = 5'ha == opcode ? retarg_5 : _GEN_518; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_557 = 5'ha == opcode ? retarg_6 : _GEN_519; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_558 = 5'ha == opcode ? retarg_7 : _GEN_520; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_559 = 5'ha == opcode ? hfutex_masks_0_0 : _GEN_521; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_560 = 5'ha == opcode ? hfutex_masks_0_1 : _GEN_522; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_561 = 5'ha == opcode ? hfutex_masks_0_2 : _GEN_523; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_562 = 5'ha == opcode ? hfutex_masks_0_3 : _GEN_524; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_563 = 5'ha == opcode ? hfutex_masks_1_0 : _GEN_525; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_564 = 5'ha == opcode ? hfutex_masks_1_1 : _GEN_526; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_565 = 5'ha == opcode ? hfutex_masks_1_2 : _GEN_527; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_566 = 5'ha == opcode ? hfutex_masks_1_3 : _GEN_528; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_567 = 5'ha == opcode ? hfutex_masks_2_0 : _GEN_529; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_568 = 5'ha == opcode ? hfutex_masks_2_1 : _GEN_530; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_569 = 5'ha == opcode ? hfutex_masks_2_2 : _GEN_531; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_570 = 5'ha == opcode ? hfutex_masks_2_3 : _GEN_532; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_571 = 5'ha == opcode ? hfutex_masks_3_0 : _GEN_533; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_572 = 5'ha == opcode ? hfutex_masks_3_1 : _GEN_534; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_573 = 5'ha == opcode ? hfutex_masks_3_2 : _GEN_535; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_574 = 5'ha == opcode ? hfutex_masks_3_3 : _GEN_536; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_575 = 5'ha == opcode ? hfutex_pos_0 : _GEN_537; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_576 = 5'ha == opcode ? hfutex_pos_1 : _GEN_538; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_577 = 5'ha == opcode ? hfutex_pos_2 : _GEN_539; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_578 = 5'ha == opcode ? hfutex_pos_3 : _GEN_540; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_579 = 5'ha == opcode ? send_hear : _GEN_541; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_580 = 5'h9 == opcode ? 5'hf : _GEN_542; // @[NulCtrlMP.scala 236:24 255:37]
  wire [7:0] _GEN_581 = 5'h9 == opcode ? _GEN_133 : _GEN_543; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_582 = 5'h9 == opcode ? _GEN_134 : _GEN_544; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_583 = 5'h9 == opcode ? _GEN_135 : _GEN_545; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_584 = 5'h9 == opcode ? _GEN_136 : _GEN_546; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_585 = 5'h9 == opcode ? _GEN_137 : _GEN_547; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_586 = 5'h9 == opcode ? _GEN_138 : _GEN_548; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_587 = 5'h9 == opcode ? _GEN_139 : _GEN_549; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_588 = 5'h9 == opcode ? _GEN_140 : _GEN_550; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_589 = 5'h9 == opcode ? retarg_0 : _GEN_551; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_590 = 5'h9 == opcode ? retarg_1 : _GEN_552; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_591 = 5'h9 == opcode ? retarg_2 : _GEN_553; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_592 = 5'h9 == opcode ? retarg_3 : _GEN_554; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_593 = 5'h9 == opcode ? retarg_4 : _GEN_555; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_594 = 5'h9 == opcode ? retarg_5 : _GEN_556; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_595 = 5'h9 == opcode ? retarg_6 : _GEN_557; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_596 = 5'h9 == opcode ? retarg_7 : _GEN_558; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_597 = 5'h9 == opcode ? hfutex_masks_0_0 : _GEN_559; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_598 = 5'h9 == opcode ? hfutex_masks_0_1 : _GEN_560; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_599 = 5'h9 == opcode ? hfutex_masks_0_2 : _GEN_561; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_600 = 5'h9 == opcode ? hfutex_masks_0_3 : _GEN_562; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_601 = 5'h9 == opcode ? hfutex_masks_1_0 : _GEN_563; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_602 = 5'h9 == opcode ? hfutex_masks_1_1 : _GEN_564; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_603 = 5'h9 == opcode ? hfutex_masks_1_2 : _GEN_565; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_604 = 5'h9 == opcode ? hfutex_masks_1_3 : _GEN_566; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_605 = 5'h9 == opcode ? hfutex_masks_2_0 : _GEN_567; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_606 = 5'h9 == opcode ? hfutex_masks_2_1 : _GEN_568; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_607 = 5'h9 == opcode ? hfutex_masks_2_2 : _GEN_569; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_608 = 5'h9 == opcode ? hfutex_masks_2_3 : _GEN_570; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_609 = 5'h9 == opcode ? hfutex_masks_3_0 : _GEN_571; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_610 = 5'h9 == opcode ? hfutex_masks_3_1 : _GEN_572; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_611 = 5'h9 == opcode ? hfutex_masks_3_2 : _GEN_573; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_612 = 5'h9 == opcode ? hfutex_masks_3_3 : _GEN_574; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_613 = 5'h9 == opcode ? hfutex_pos_0 : _GEN_575; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_614 = 5'h9 == opcode ? hfutex_pos_1 : _GEN_576; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_615 = 5'h9 == opcode ? hfutex_pos_2 : _GEN_577; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_616 = 5'h9 == opcode ? hfutex_pos_3 : _GEN_578; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_617 = 5'h9 == opcode ? send_hear : _GEN_579; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_618 = 5'h8 == opcode ? 5'he : _GEN_580; // @[NulCtrlMP.scala 236:24 254:37]
  wire [7:0] _GEN_619 = 5'h8 == opcode ? _GEN_133 : _GEN_581; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_620 = 5'h8 == opcode ? _GEN_134 : _GEN_582; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_621 = 5'h8 == opcode ? _GEN_135 : _GEN_583; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_622 = 5'h8 == opcode ? _GEN_136 : _GEN_584; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_623 = 5'h8 == opcode ? _GEN_137 : _GEN_585; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_624 = 5'h8 == opcode ? _GEN_138 : _GEN_586; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_625 = 5'h8 == opcode ? _GEN_139 : _GEN_587; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_626 = 5'h8 == opcode ? _GEN_140 : _GEN_588; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_627 = 5'h8 == opcode ? retarg_0 : _GEN_589; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_628 = 5'h8 == opcode ? retarg_1 : _GEN_590; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_629 = 5'h8 == opcode ? retarg_2 : _GEN_591; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_630 = 5'h8 == opcode ? retarg_3 : _GEN_592; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_631 = 5'h8 == opcode ? retarg_4 : _GEN_593; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_632 = 5'h8 == opcode ? retarg_5 : _GEN_594; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_633 = 5'h8 == opcode ? retarg_6 : _GEN_595; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_634 = 5'h8 == opcode ? retarg_7 : _GEN_596; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_635 = 5'h8 == opcode ? hfutex_masks_0_0 : _GEN_597; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_636 = 5'h8 == opcode ? hfutex_masks_0_1 : _GEN_598; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_637 = 5'h8 == opcode ? hfutex_masks_0_2 : _GEN_599; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_638 = 5'h8 == opcode ? hfutex_masks_0_3 : _GEN_600; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_639 = 5'h8 == opcode ? hfutex_masks_1_0 : _GEN_601; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_640 = 5'h8 == opcode ? hfutex_masks_1_1 : _GEN_602; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_641 = 5'h8 == opcode ? hfutex_masks_1_2 : _GEN_603; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_642 = 5'h8 == opcode ? hfutex_masks_1_3 : _GEN_604; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_643 = 5'h8 == opcode ? hfutex_masks_2_0 : _GEN_605; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_644 = 5'h8 == opcode ? hfutex_masks_2_1 : _GEN_606; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_645 = 5'h8 == opcode ? hfutex_masks_2_2 : _GEN_607; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_646 = 5'h8 == opcode ? hfutex_masks_2_3 : _GEN_608; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_647 = 5'h8 == opcode ? hfutex_masks_3_0 : _GEN_609; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_648 = 5'h8 == opcode ? hfutex_masks_3_1 : _GEN_610; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_649 = 5'h8 == opcode ? hfutex_masks_3_2 : _GEN_611; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_650 = 5'h8 == opcode ? hfutex_masks_3_3 : _GEN_612; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_651 = 5'h8 == opcode ? hfutex_pos_0 : _GEN_613; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_652 = 5'h8 == opcode ? hfutex_pos_1 : _GEN_614; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_653 = 5'h8 == opcode ? hfutex_pos_2 : _GEN_615; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_654 = 5'h8 == opcode ? hfutex_pos_3 : _GEN_616; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_655 = 5'h8 == opcode ? send_hear : _GEN_617; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_656 = 5'h7 == opcode ? 5'h16 : _GEN_618; // @[NulCtrlMP.scala 236:24 253:37]
  wire [7:0] _GEN_657 = 5'h7 == opcode ? _GEN_133 : _GEN_619; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_658 = 5'h7 == opcode ? _GEN_134 : _GEN_620; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_659 = 5'h7 == opcode ? _GEN_135 : _GEN_621; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_660 = 5'h7 == opcode ? _GEN_136 : _GEN_622; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_661 = 5'h7 == opcode ? _GEN_137 : _GEN_623; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_662 = 5'h7 == opcode ? _GEN_138 : _GEN_624; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_663 = 5'h7 == opcode ? _GEN_139 : _GEN_625; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_664 = 5'h7 == opcode ? _GEN_140 : _GEN_626; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_665 = 5'h7 == opcode ? retarg_0 : _GEN_627; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_666 = 5'h7 == opcode ? retarg_1 : _GEN_628; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_667 = 5'h7 == opcode ? retarg_2 : _GEN_629; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_668 = 5'h7 == opcode ? retarg_3 : _GEN_630; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_669 = 5'h7 == opcode ? retarg_4 : _GEN_631; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_670 = 5'h7 == opcode ? retarg_5 : _GEN_632; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_671 = 5'h7 == opcode ? retarg_6 : _GEN_633; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_672 = 5'h7 == opcode ? retarg_7 : _GEN_634; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_673 = 5'h7 == opcode ? hfutex_masks_0_0 : _GEN_635; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_674 = 5'h7 == opcode ? hfutex_masks_0_1 : _GEN_636; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_675 = 5'h7 == opcode ? hfutex_masks_0_2 : _GEN_637; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_676 = 5'h7 == opcode ? hfutex_masks_0_3 : _GEN_638; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_677 = 5'h7 == opcode ? hfutex_masks_1_0 : _GEN_639; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_678 = 5'h7 == opcode ? hfutex_masks_1_1 : _GEN_640; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_679 = 5'h7 == opcode ? hfutex_masks_1_2 : _GEN_641; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_680 = 5'h7 == opcode ? hfutex_masks_1_3 : _GEN_642; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_681 = 5'h7 == opcode ? hfutex_masks_2_0 : _GEN_643; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_682 = 5'h7 == opcode ? hfutex_masks_2_1 : _GEN_644; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_683 = 5'h7 == opcode ? hfutex_masks_2_2 : _GEN_645; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_684 = 5'h7 == opcode ? hfutex_masks_2_3 : _GEN_646; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_685 = 5'h7 == opcode ? hfutex_masks_3_0 : _GEN_647; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_686 = 5'h7 == opcode ? hfutex_masks_3_1 : _GEN_648; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_687 = 5'h7 == opcode ? hfutex_masks_3_2 : _GEN_649; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_688 = 5'h7 == opcode ? hfutex_masks_3_3 : _GEN_650; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_689 = 5'h7 == opcode ? hfutex_pos_0 : _GEN_651; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_690 = 5'h7 == opcode ? hfutex_pos_1 : _GEN_652; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_691 = 5'h7 == opcode ? hfutex_pos_2 : _GEN_653; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_692 = 5'h7 == opcode ? hfutex_pos_3 : _GEN_654; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_693 = 5'h7 == opcode ? send_hear : _GEN_655; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_694 = 5'h6 == opcode ? 5'hd : _GEN_656; // @[NulCtrlMP.scala 236:24 252:37]
  wire [7:0] _GEN_695 = 5'h6 == opcode ? _GEN_133 : _GEN_657; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_696 = 5'h6 == opcode ? _GEN_134 : _GEN_658; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_697 = 5'h6 == opcode ? _GEN_135 : _GEN_659; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_698 = 5'h6 == opcode ? _GEN_136 : _GEN_660; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_699 = 5'h6 == opcode ? _GEN_137 : _GEN_661; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_700 = 5'h6 == opcode ? _GEN_138 : _GEN_662; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_701 = 5'h6 == opcode ? _GEN_139 : _GEN_663; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_702 = 5'h6 == opcode ? _GEN_140 : _GEN_664; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_703 = 5'h6 == opcode ? retarg_0 : _GEN_665; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_704 = 5'h6 == opcode ? retarg_1 : _GEN_666; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_705 = 5'h6 == opcode ? retarg_2 : _GEN_667; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_706 = 5'h6 == opcode ? retarg_3 : _GEN_668; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_707 = 5'h6 == opcode ? retarg_4 : _GEN_669; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_708 = 5'h6 == opcode ? retarg_5 : _GEN_670; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_709 = 5'h6 == opcode ? retarg_6 : _GEN_671; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_710 = 5'h6 == opcode ? retarg_7 : _GEN_672; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_711 = 5'h6 == opcode ? hfutex_masks_0_0 : _GEN_673; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_712 = 5'h6 == opcode ? hfutex_masks_0_1 : _GEN_674; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_713 = 5'h6 == opcode ? hfutex_masks_0_2 : _GEN_675; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_714 = 5'h6 == opcode ? hfutex_masks_0_3 : _GEN_676; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_715 = 5'h6 == opcode ? hfutex_masks_1_0 : _GEN_677; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_716 = 5'h6 == opcode ? hfutex_masks_1_1 : _GEN_678; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_717 = 5'h6 == opcode ? hfutex_masks_1_2 : _GEN_679; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_718 = 5'h6 == opcode ? hfutex_masks_1_3 : _GEN_680; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_719 = 5'h6 == opcode ? hfutex_masks_2_0 : _GEN_681; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_720 = 5'h6 == opcode ? hfutex_masks_2_1 : _GEN_682; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_721 = 5'h6 == opcode ? hfutex_masks_2_2 : _GEN_683; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_722 = 5'h6 == opcode ? hfutex_masks_2_3 : _GEN_684; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_723 = 5'h6 == opcode ? hfutex_masks_3_0 : _GEN_685; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_724 = 5'h6 == opcode ? hfutex_masks_3_1 : _GEN_686; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_725 = 5'h6 == opcode ? hfutex_masks_3_2 : _GEN_687; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_726 = 5'h6 == opcode ? hfutex_masks_3_3 : _GEN_688; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_727 = 5'h6 == opcode ? hfutex_pos_0 : _GEN_689; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_728 = 5'h6 == opcode ? hfutex_pos_1 : _GEN_690; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_729 = 5'h6 == opcode ? hfutex_pos_2 : _GEN_691; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_730 = 5'h6 == opcode ? hfutex_pos_3 : _GEN_692; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_731 = 5'h6 == opcode ? send_hear : _GEN_693; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_732 = 5'h5 == opcode ? 5'hc : _GEN_694; // @[NulCtrlMP.scala 236:24 251:36]
  wire [7:0] _GEN_733 = 5'h5 == opcode ? _GEN_133 : _GEN_695; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_734 = 5'h5 == opcode ? _GEN_134 : _GEN_696; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_735 = 5'h5 == opcode ? _GEN_135 : _GEN_697; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_736 = 5'h5 == opcode ? _GEN_136 : _GEN_698; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_737 = 5'h5 == opcode ? _GEN_137 : _GEN_699; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_738 = 5'h5 == opcode ? _GEN_138 : _GEN_700; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_739 = 5'h5 == opcode ? _GEN_139 : _GEN_701; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_740 = 5'h5 == opcode ? _GEN_140 : _GEN_702; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_741 = 5'h5 == opcode ? retarg_0 : _GEN_703; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_742 = 5'h5 == opcode ? retarg_1 : _GEN_704; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_743 = 5'h5 == opcode ? retarg_2 : _GEN_705; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_744 = 5'h5 == opcode ? retarg_3 : _GEN_706; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_745 = 5'h5 == opcode ? retarg_4 : _GEN_707; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_746 = 5'h5 == opcode ? retarg_5 : _GEN_708; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_747 = 5'h5 == opcode ? retarg_6 : _GEN_709; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_748 = 5'h5 == opcode ? retarg_7 : _GEN_710; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_749 = 5'h5 == opcode ? hfutex_masks_0_0 : _GEN_711; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_750 = 5'h5 == opcode ? hfutex_masks_0_1 : _GEN_712; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_751 = 5'h5 == opcode ? hfutex_masks_0_2 : _GEN_713; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_752 = 5'h5 == opcode ? hfutex_masks_0_3 : _GEN_714; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_753 = 5'h5 == opcode ? hfutex_masks_1_0 : _GEN_715; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_754 = 5'h5 == opcode ? hfutex_masks_1_1 : _GEN_716; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_755 = 5'h5 == opcode ? hfutex_masks_1_2 : _GEN_717; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_756 = 5'h5 == opcode ? hfutex_masks_1_3 : _GEN_718; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_757 = 5'h5 == opcode ? hfutex_masks_2_0 : _GEN_719; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_758 = 5'h5 == opcode ? hfutex_masks_2_1 : _GEN_720; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_759 = 5'h5 == opcode ? hfutex_masks_2_2 : _GEN_721; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_760 = 5'h5 == opcode ? hfutex_masks_2_3 : _GEN_722; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_761 = 5'h5 == opcode ? hfutex_masks_3_0 : _GEN_723; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_762 = 5'h5 == opcode ? hfutex_masks_3_1 : _GEN_724; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_763 = 5'h5 == opcode ? hfutex_masks_3_2 : _GEN_725; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_764 = 5'h5 == opcode ? hfutex_masks_3_3 : _GEN_726; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_765 = 5'h5 == opcode ? hfutex_pos_0 : _GEN_727; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_766 = 5'h5 == opcode ? hfutex_pos_1 : _GEN_728; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_767 = 5'h5 == opcode ? hfutex_pos_2 : _GEN_729; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_768 = 5'h5 == opcode ? hfutex_pos_3 : _GEN_730; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_769 = 5'h5 == opcode ? send_hear : _GEN_731; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_770 = 5'h4 == opcode ? {{1'd0}, _GEN_161} : _GEN_732; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_771 = 5'h4 == opcode ? _GEN_133 : _GEN_733; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_772 = 5'h4 == opcode ? _GEN_134 : _GEN_734; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_773 = 5'h4 == opcode ? _GEN_135 : _GEN_735; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_774 = 5'h4 == opcode ? _GEN_136 : _GEN_736; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_775 = 5'h4 == opcode ? _GEN_137 : _GEN_737; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_776 = 5'h4 == opcode ? _GEN_138 : _GEN_738; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_777 = 5'h4 == opcode ? _GEN_139 : _GEN_739; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_778 = 5'h4 == opcode ? _GEN_140 : _GEN_740; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_779 = 5'h4 == opcode ? retarg_0 : _GEN_741; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_780 = 5'h4 == opcode ? retarg_1 : _GEN_742; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_781 = 5'h4 == opcode ? retarg_2 : _GEN_743; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_782 = 5'h4 == opcode ? retarg_3 : _GEN_744; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_783 = 5'h4 == opcode ? retarg_4 : _GEN_745; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_784 = 5'h4 == opcode ? retarg_5 : _GEN_746; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_785 = 5'h4 == opcode ? retarg_6 : _GEN_747; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_786 = 5'h4 == opcode ? retarg_7 : _GEN_748; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_787 = 5'h4 == opcode ? hfutex_masks_0_0 : _GEN_749; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_788 = 5'h4 == opcode ? hfutex_masks_0_1 : _GEN_750; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_789 = 5'h4 == opcode ? hfutex_masks_0_2 : _GEN_751; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_790 = 5'h4 == opcode ? hfutex_masks_0_3 : _GEN_752; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_791 = 5'h4 == opcode ? hfutex_masks_1_0 : _GEN_753; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_792 = 5'h4 == opcode ? hfutex_masks_1_1 : _GEN_754; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_793 = 5'h4 == opcode ? hfutex_masks_1_2 : _GEN_755; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_794 = 5'h4 == opcode ? hfutex_masks_1_3 : _GEN_756; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_795 = 5'h4 == opcode ? hfutex_masks_2_0 : _GEN_757; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_796 = 5'h4 == opcode ? hfutex_masks_2_1 : _GEN_758; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_797 = 5'h4 == opcode ? hfutex_masks_2_2 : _GEN_759; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_798 = 5'h4 == opcode ? hfutex_masks_2_3 : _GEN_760; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_799 = 5'h4 == opcode ? hfutex_masks_3_0 : _GEN_761; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_800 = 5'h4 == opcode ? hfutex_masks_3_1 : _GEN_762; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_801 = 5'h4 == opcode ? hfutex_masks_3_2 : _GEN_763; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_802 = 5'h4 == opcode ? hfutex_masks_3_3 : _GEN_764; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_803 = 5'h4 == opcode ? hfutex_pos_0 : _GEN_765; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_804 = 5'h4 == opcode ? hfutex_pos_1 : _GEN_766; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_805 = 5'h4 == opcode ? hfutex_pos_2 : _GEN_767; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_806 = 5'h4 == opcode ? hfutex_pos_3 : _GEN_768; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_807 = 5'h4 == opcode ? send_hear : _GEN_769; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_808 = 5'h3 == opcode ? 5'ha : _GEN_770; // @[NulCtrlMP.scala 236:24 245:35]
  wire [7:0] _GEN_809 = 5'h3 == opcode ? _GEN_133 : _GEN_771; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_810 = 5'h3 == opcode ? _GEN_134 : _GEN_772; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_811 = 5'h3 == opcode ? _GEN_135 : _GEN_773; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_812 = 5'h3 == opcode ? _GEN_136 : _GEN_774; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_813 = 5'h3 == opcode ? _GEN_137 : _GEN_775; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_814 = 5'h3 == opcode ? _GEN_138 : _GEN_776; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_815 = 5'h3 == opcode ? _GEN_139 : _GEN_777; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_816 = 5'h3 == opcode ? _GEN_140 : _GEN_778; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_817 = 5'h3 == opcode ? retarg_0 : _GEN_779; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_818 = 5'h3 == opcode ? retarg_1 : _GEN_780; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_819 = 5'h3 == opcode ? retarg_2 : _GEN_781; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_820 = 5'h3 == opcode ? retarg_3 : _GEN_782; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_821 = 5'h3 == opcode ? retarg_4 : _GEN_783; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_822 = 5'h3 == opcode ? retarg_5 : _GEN_784; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_823 = 5'h3 == opcode ? retarg_6 : _GEN_785; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_824 = 5'h3 == opcode ? retarg_7 : _GEN_786; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_825 = 5'h3 == opcode ? hfutex_masks_0_0 : _GEN_787; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_826 = 5'h3 == opcode ? hfutex_masks_0_1 : _GEN_788; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_827 = 5'h3 == opcode ? hfutex_masks_0_2 : _GEN_789; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_828 = 5'h3 == opcode ? hfutex_masks_0_3 : _GEN_790; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_829 = 5'h3 == opcode ? hfutex_masks_1_0 : _GEN_791; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_830 = 5'h3 == opcode ? hfutex_masks_1_1 : _GEN_792; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_831 = 5'h3 == opcode ? hfutex_masks_1_2 : _GEN_793; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_832 = 5'h3 == opcode ? hfutex_masks_1_3 : _GEN_794; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_833 = 5'h3 == opcode ? hfutex_masks_2_0 : _GEN_795; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_834 = 5'h3 == opcode ? hfutex_masks_2_1 : _GEN_796; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_835 = 5'h3 == opcode ? hfutex_masks_2_2 : _GEN_797; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_836 = 5'h3 == opcode ? hfutex_masks_2_3 : _GEN_798; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_837 = 5'h3 == opcode ? hfutex_masks_3_0 : _GEN_799; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_838 = 5'h3 == opcode ? hfutex_masks_3_1 : _GEN_800; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_839 = 5'h3 == opcode ? hfutex_masks_3_2 : _GEN_801; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_840 = 5'h3 == opcode ? hfutex_masks_3_3 : _GEN_802; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_841 = 5'h3 == opcode ? hfutex_pos_0 : _GEN_803; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_842 = 5'h3 == opcode ? hfutex_pos_1 : _GEN_804; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_843 = 5'h3 == opcode ? hfutex_pos_2 : _GEN_805; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_844 = 5'h3 == opcode ? hfutex_pos_3 : _GEN_806; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_845 = 5'h3 == opcode ? send_hear : _GEN_807; // @[NulCtrlMP.scala 236:24 169:28]
  wire  _GEN_846 = 5'h2 == opcode & _GEN_145; // @[NulCtrlMP.scala 236:24 44:27]
  wire  _GEN_847 = 5'h2 == opcode & _GEN_146; // @[NulCtrlMP.scala 236:24 44:27]
  wire  _GEN_848 = 5'h2 == opcode & _GEN_147; // @[NulCtrlMP.scala 236:24 44:27]
  wire  _GEN_849 = 5'h2 == opcode & _GEN_148; // @[NulCtrlMP.scala 236:24 44:27]
  wire [4:0] _GEN_850 = 5'h2 == opcode ? 5'h5 : _GEN_808; // @[NulCtrlMP.scala 235:15 236:24]
  wire [7:0] _GEN_851 = 5'h2 == opcode ? _GEN_133 : _GEN_809; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_852 = 5'h2 == opcode ? _GEN_134 : _GEN_810; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_853 = 5'h2 == opcode ? _GEN_135 : _GEN_811; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_854 = 5'h2 == opcode ? _GEN_136 : _GEN_812; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_855 = 5'h2 == opcode ? _GEN_137 : _GEN_813; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_856 = 5'h2 == opcode ? _GEN_138 : _GEN_814; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_857 = 5'h2 == opcode ? _GEN_139 : _GEN_815; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_858 = 5'h2 == opcode ? _GEN_140 : _GEN_816; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_859 = 5'h2 == opcode ? retarg_0 : _GEN_817; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_860 = 5'h2 == opcode ? retarg_1 : _GEN_818; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_861 = 5'h2 == opcode ? retarg_2 : _GEN_819; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_862 = 5'h2 == opcode ? retarg_3 : _GEN_820; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_863 = 5'h2 == opcode ? retarg_4 : _GEN_821; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_864 = 5'h2 == opcode ? retarg_5 : _GEN_822; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_865 = 5'h2 == opcode ? retarg_6 : _GEN_823; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_866 = 5'h2 == opcode ? retarg_7 : _GEN_824; // @[NulCtrlMP.scala 236:24 152:25]
  wire [47:0] _GEN_867 = 5'h2 == opcode ? hfutex_masks_0_0 : _GEN_825; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_868 = 5'h2 == opcode ? hfutex_masks_0_1 : _GEN_826; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_869 = 5'h2 == opcode ? hfutex_masks_0_2 : _GEN_827; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_870 = 5'h2 == opcode ? hfutex_masks_0_3 : _GEN_828; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_871 = 5'h2 == opcode ? hfutex_masks_1_0 : _GEN_829; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_872 = 5'h2 == opcode ? hfutex_masks_1_1 : _GEN_830; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_873 = 5'h2 == opcode ? hfutex_masks_1_2 : _GEN_831; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_874 = 5'h2 == opcode ? hfutex_masks_1_3 : _GEN_832; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_875 = 5'h2 == opcode ? hfutex_masks_2_0 : _GEN_833; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_876 = 5'h2 == opcode ? hfutex_masks_2_1 : _GEN_834; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_877 = 5'h2 == opcode ? hfutex_masks_2_2 : _GEN_835; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_878 = 5'h2 == opcode ? hfutex_masks_2_3 : _GEN_836; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_879 = 5'h2 == opcode ? hfutex_masks_3_0 : _GEN_837; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_880 = 5'h2 == opcode ? hfutex_masks_3_1 : _GEN_838; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_881 = 5'h2 == opcode ? hfutex_masks_3_2 : _GEN_839; // @[NulCtrlMP.scala 236:24 162:31]
  wire [47:0] _GEN_882 = 5'h2 == opcode ? hfutex_masks_3_3 : _GEN_840; // @[NulCtrlMP.scala 236:24 162:31]
  wire [1:0] _GEN_883 = 5'h2 == opcode ? hfutex_pos_0 : _GEN_841; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_884 = 5'h2 == opcode ? hfutex_pos_1 : _GEN_842; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_885 = 5'h2 == opcode ? hfutex_pos_2 : _GEN_843; // @[NulCtrlMP.scala 236:24 163:29]
  wire [1:0] _GEN_886 = 5'h2 == opcode ? hfutex_pos_3 : _GEN_844; // @[NulCtrlMP.scala 236:24 163:29]
  wire  _GEN_887 = 5'h2 == opcode ? send_hear : _GEN_845; // @[NulCtrlMP.scala 236:24 169:28]
  wire  _GEN_888 = 5'h1 == opcode ? _GEN_145 : _GEN_846; // @[NulCtrlMP.scala 236:24]
  wire  _GEN_889 = 5'h1 == opcode ? _GEN_146 : _GEN_847; // @[NulCtrlMP.scala 236:24]
  wire  _GEN_890 = 5'h1 == opcode ? _GEN_147 : _GEN_848; // @[NulCtrlMP.scala 236:24]
  wire  _GEN_891 = 5'h1 == opcode ? _GEN_148 : _GEN_849; // @[NulCtrlMP.scala 236:24]
  wire [1:0] _GEN_892 = 5'h1 == opcode ? _GEN_149 : _GEN_21; // @[NulCtrlMP.scala 236:24]
  wire [1:0] _GEN_893 = 5'h1 == opcode ? _GEN_150 : _GEN_22; // @[NulCtrlMP.scala 236:24]
  wire [1:0] _GEN_894 = 5'h1 == opcode ? _GEN_151 : _GEN_23; // @[NulCtrlMP.scala 236:24]
  wire [1:0] _GEN_895 = 5'h1 == opcode ? _GEN_152 : _GEN_24; // @[NulCtrlMP.scala 236:24]
  wire [4:0] _GEN_896 = 5'h1 == opcode ? 5'h5 : _GEN_850; // @[NulCtrlMP.scala 235:15 236:24]
  wire [7:0] _GEN_905 = 5'h1 == opcode ? retarg_0 : _GEN_859; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_906 = 5'h1 == opcode ? retarg_1 : _GEN_860; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_907 = 5'h1 == opcode ? retarg_2 : _GEN_861; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_908 = 5'h1 == opcode ? retarg_3 : _GEN_862; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_909 = 5'h1 == opcode ? retarg_4 : _GEN_863; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_910 = 5'h1 == opcode ? retarg_5 : _GEN_864; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_911 = 5'h1 == opcode ? retarg_6 : _GEN_865; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_912 = 5'h1 == opcode ? retarg_7 : _GEN_866; // @[NulCtrlMP.scala 236:24 152:25]
  wire  _GEN_933 = 5'h1 == opcode ? send_hear : _GEN_887; // @[NulCtrlMP.scala 236:24 169:28]
  wire [4:0] _GEN_934 = 5'h0 == opcode ? 5'h8 : _GEN_896; // @[NulCtrlMP.scala 236:24 237:36]
  wire  _GEN_935 = 5'h0 == opcode ? 1'h0 : _GEN_888; // @[NulCtrlMP.scala 236:24 44:27]
  wire  _GEN_936 = 5'h0 == opcode ? 1'h0 : _GEN_889; // @[NulCtrlMP.scala 236:24 44:27]
  wire  _GEN_937 = 5'h0 == opcode ? 1'h0 : _GEN_890; // @[NulCtrlMP.scala 236:24 44:27]
  wire  _GEN_938 = 5'h0 == opcode ? 1'h0 : _GEN_891; // @[NulCtrlMP.scala 236:24 44:27]
  wire [1:0] _GEN_939 = 5'h0 == opcode ? _GEN_21 : _GEN_892; // @[NulCtrlMP.scala 236:24]
  wire [1:0] _GEN_940 = 5'h0 == opcode ? _GEN_22 : _GEN_893; // @[NulCtrlMP.scala 236:24]
  wire [1:0] _GEN_941 = 5'h0 == opcode ? _GEN_23 : _GEN_894; // @[NulCtrlMP.scala 236:24]
  wire [1:0] _GEN_942 = 5'h0 == opcode ? _GEN_24 : _GEN_895; // @[NulCtrlMP.scala 236:24]
  wire [7:0] _GEN_951 = 5'h0 == opcode ? retarg_0 : _GEN_905; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_952 = 5'h0 == opcode ? retarg_1 : _GEN_906; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_953 = 5'h0 == opcode ? retarg_2 : _GEN_907; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_954 = 5'h0 == opcode ? retarg_3 : _GEN_908; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_955 = 5'h0 == opcode ? retarg_4 : _GEN_909; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_956 = 5'h0 == opcode ? retarg_5 : _GEN_910; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_957 = 5'h0 == opcode ? retarg_6 : _GEN_911; // @[NulCtrlMP.scala 236:24 152:25]
  wire [7:0] _GEN_958 = 5'h0 == opcode ? retarg_7 : _GEN_912; // @[NulCtrlMP.scala 236:24 152:25]
  wire  _GEN_979 = 5'h0 == opcode ? send_hear : _GEN_933; // @[NulCtrlMP.scala 236:24 169:28]
  wire [7:0] _GEN_981 = 4'h1 == trans_pos[3:0] ? io_rx_bits : _GEN_127; // @[NulCtrlMP.scala 296:{26,26}]
  wire [7:0] _GEN_997 = _T_66 & io_rx_valid ? _GEN_981 : _GEN_127; // @[NulCtrlMP.scala 295:57]
  wire [9:0] _GEN_1012 = _T_66 & io_rx_valid ? _T_69 : _GEN_142; // @[NulCtrlMP.scala 295:57 297:19]
  wire [9:0] _GEN_1013 = state == 5'h4 ? 10'h1 : _GEN_143; // @[NulCtrlMP.scala 232:33 233:21]
  wire [9:0] _GEN_1014 = state == 5'h4 ? 10'h1 : _GEN_1012; // @[NulCtrlMP.scala 232:33 234:19]
  wire [4:0] _GEN_1015 = state == 5'h4 ? _GEN_934 : _GEN_144; // @[NulCtrlMP.scala 232:33]
  wire [1:0] _GEN_1020 = state == 5'h4 ? _GEN_939 : _GEN_21; // @[NulCtrlMP.scala 232:33]
  wire [1:0] _GEN_1021 = state == 5'h4 ? _GEN_940 : _GEN_22; // @[NulCtrlMP.scala 232:33]
  wire [1:0] _GEN_1022 = state == 5'h4 ? _GEN_941 : _GEN_23; // @[NulCtrlMP.scala 232:33]
  wire [1:0] _GEN_1023 = state == 5'h4 ? _GEN_942 : _GEN_24; // @[NulCtrlMP.scala 232:33]
  wire [7:0] _GEN_1032 = state == 5'h4 ? _GEN_951 : retarg_0; // @[NulCtrlMP.scala 152:25 232:33]
  wire [7:0] _GEN_1033 = state == 5'h4 ? _GEN_952 : retarg_1; // @[NulCtrlMP.scala 152:25 232:33]
  wire [7:0] _GEN_1034 = state == 5'h4 ? _GEN_953 : retarg_2; // @[NulCtrlMP.scala 152:25 232:33]
  wire [7:0] _GEN_1035 = state == 5'h4 ? _GEN_954 : retarg_3; // @[NulCtrlMP.scala 152:25 232:33]
  wire [7:0] _GEN_1036 = state == 5'h4 ? _GEN_955 : retarg_4; // @[NulCtrlMP.scala 152:25 232:33]
  wire [7:0] _GEN_1037 = state == 5'h4 ? _GEN_956 : retarg_5; // @[NulCtrlMP.scala 152:25 232:33]
  wire [7:0] _GEN_1038 = state == 5'h4 ? _GEN_957 : retarg_6; // @[NulCtrlMP.scala 152:25 232:33]
  wire [7:0] _GEN_1039 = state == 5'h4 ? _GEN_958 : retarg_7; // @[NulCtrlMP.scala 152:25 232:33]
  wire  _GEN_1060 = state == 5'h4 ? _GEN_979 : send_hear; // @[NulCtrlMP.scala 169:28 232:33]
  wire [7:0] _GEN_1062 = state == 5'h4 ? _GEN_127 : _GEN_997; // @[NulCtrlMP.scala 232:33]
  wire  _T_102 = state == 5'h5; // @[NulCtrlMP.scala 300:16]
  wire [7:0] _io_tx_bits_T = {opoff,opcode}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_1069 = opcode == 5'h8 | opcode == 5'ha | opcode == 5'h10 | opcode == 5'h11 ? 4'h8 : 4'h0; // @[NulCtrlMP.scala 308:123 309:29 312:29]
  wire [4:0] _GEN_1070 = opcode == 5'h8 | opcode == 5'ha | opcode == 5'h10 | opcode == 5'h11 ? 5'h6 : 5'h1f; // @[NulCtrlMP.scala 308:123 310:23 313:23]
  wire [3:0] _GEN_1071 = opcode == 5'h0 ? 4'he : _GEN_1069; // @[NulCtrlMP.scala 305:41 306:29]
  wire [4:0] _GEN_1072 = opcode == 5'h0 ? 5'h6 : _GEN_1070; // @[NulCtrlMP.scala 305:41 307:23]
  wire [9:0] _GEN_1073 = io_tx_ready ? {{6'd0}, _GEN_1071} : _GEN_1013; // @[NulCtrlMP.scala 304:27]
  wire [4:0] _GEN_1074 = io_tx_ready ? _GEN_1072 : _GEN_1015; // @[NulCtrlMP.scala 304:27]
  wire [7:0] _GEN_1076 = state == 5'h5 ? _io_tx_bits_T : 8'h0; // @[NulCtrlMP.scala 300:37 302:20 34:16]
  wire [9:0] _GEN_1077 = state == 5'h5 ? 10'h0 : _GEN_1014; // @[NulCtrlMP.scala 300:37 303:19]
  wire [9:0] _GEN_1078 = state == 5'h5 ? _GEN_1073 : _GEN_1013; // @[NulCtrlMP.scala 300:37]
  wire [4:0] _GEN_1079 = state == 5'h5 ? _GEN_1074 : _GEN_1015; // @[NulCtrlMP.scala 300:37]
  wire [7:0] _GEN_1081 = 4'h1 == trans_pos[3:0] ? retarg_1 : retarg_0; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1082 = 4'h2 == trans_pos[3:0] ? retarg_2 : _GEN_1081; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1083 = 4'h3 == trans_pos[3:0] ? retarg_3 : _GEN_1082; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1084 = 4'h4 == trans_pos[3:0] ? retarg_4 : _GEN_1083; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1085 = 4'h5 == trans_pos[3:0] ? retarg_5 : _GEN_1084; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1086 = 4'h6 == trans_pos[3:0] ? retarg_6 : _GEN_1085; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1087 = 4'h7 == trans_pos[3:0] ? retarg_7 : _GEN_1086; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1088 = 4'h8 == trans_pos[3:0] ? retarg_8 : _GEN_1087; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1089 = 4'h9 == trans_pos[3:0] ? retarg_9 : _GEN_1088; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1090 = 4'ha == trans_pos[3:0] ? retarg_10 : _GEN_1089; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1091 = 4'hb == trans_pos[3:0] ? retarg_11 : _GEN_1090; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1092 = 4'hc == trans_pos[3:0] ? retarg_12 : _GEN_1091; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1093 = 4'hd == trans_pos[3:0] ? retarg_13 : _GEN_1092; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1094 = 4'he == trans_pos[3:0] ? 8'h0 : _GEN_1093; // @[NulCtrlMP.scala 320:{20,20}]
  wire [7:0] _GEN_1095 = 4'hf == trans_pos[3:0] ? 8'h0 : _GEN_1094; // @[NulCtrlMP.scala 320:{20,20}]
  wire [4:0] _GEN_1098 = _T_70 ? 5'h1f : _GEN_1079; // @[NulCtrlMP.scala 322:51 325:23]
  wire [4:0] _GEN_1101 = io_tx_ready ? _GEN_1098 : _GEN_1079; // @[NulCtrlMP.scala 321:27]
  wire  _GEN_1102 = state == 5'h6 | _T_102; // @[NulCtrlMP.scala 318:36 319:21]
  wire [7:0] _GEN_1103 = state == 5'h6 ? _GEN_1095 : _GEN_1076; // @[NulCtrlMP.scala 318:36 320:20]
  wire [4:0] _GEN_1106 = state == 5'h6 ? _GEN_1101 : _GEN_1079; // @[NulCtrlMP.scala 318:36]
  wire  all_halted = _io_cpu_0_stop_fetch_T_1 & _io_cpu_1_stop_fetch_T_1 & _io_cpu_2_stop_fetch_T_1 &
    _io_cpu_3_stop_fetch_T_1; // @[NulCtrlMP.scala 332:38]
  wire  _event_queue_io_deq_ready_T = state == 5'h8; // @[NulCtrlMP.scala 334:40]
  wire [7:0] pending_next_idx = {{6'd0}, event_queue_io_deq_bits}; // @[NulCtrlMP.scala 336:59]
  wire [7:0] _GEN_1107 = _event_queue_io_deq_ready_T & all_halted ? 8'hff : _GEN_1032; // @[NulCtrlMP.scala 340:57 341:19]
  wire [4:0] _GEN_1108 = _event_queue_io_deq_ready_T & all_halted ? 5'h5 : _GEN_1106; // @[NulCtrlMP.scala 340:57 342:15]
  wire [7:0] _GEN_1109 = _event_queue_io_deq_ready_T & event_queue_io_deq_valid ? pending_next_idx : _GEN_1062; // @[NulCtrlMP.scala 335:65 337:18]
  wire [7:0] _GEN_1110 = _event_queue_io_deq_ready_T & event_queue_io_deq_valid ? pending_next_idx : _GEN_1107; // @[NulCtrlMP.scala 335:65 338:19]
  wire [4:0] _GEN_1111 = _event_queue_io_deq_ready_T & event_queue_io_deq_valid ? 5'h9 : _GEN_1108; // @[NulCtrlMP.scala 335:65 339:15]
  reg [127:0] cnt; // @[NulCtrlMP.scala 345:22]
  reg [63:0] regback_0; // @[NulCtrlMP.scala 346:26]
  reg [63:0] regback_1; // @[NulCtrlMP.scala 346:26]
  reg [63:0] regback_2; // @[NulCtrlMP.scala 346:26]
  reg [63:0] regback_3; // @[NulCtrlMP.scala 346:26]
  reg [63:0] regback_4; // @[NulCtrlMP.scala 346:26]
  reg [63:0] regback_5; // @[NulCtrlMP.scala 346:26]
  reg [63:0] regback_6; // @[NulCtrlMP.scala 346:26]
  reg [63:0] regback_7; // @[NulCtrlMP.scala 346:26]
  reg [63:0] regback_8; // @[NulCtrlMP.scala 346:26]
  reg [63:0] regback_9; // @[NulCtrlMP.scala 346:26]
  reg [1:0] init_cnt; // @[NulCtrlMP.scala 420:27]
  wire [128:0] _cnt_T = {cnt, 1'h0}; // @[NulCtrlMP.scala 422:36]
  wire [128:0] _GEN_1112 = cnt[0] ? _cnt_T : {{1'd0}, cnt}; // @[NulCtrlMP.scala 345:22 422:{22,28}]
  wire [4:0] _GEN_1117 = 2'h0 == opidx ? 5'h7 : 5'h0; // @[NulCtrlMP.scala 370:{28,28} 47:30]
  wire [4:0] _GEN_1118 = 2'h1 == opidx ? 5'h7 : 5'h0; // @[NulCtrlMP.scala 370:{28,28} 47:30]
  wire [4:0] _GEN_1119 = 2'h2 == opidx ? 5'h7 : 5'h0; // @[NulCtrlMP.scala 370:{28,28} 47:30]
  wire [4:0] _GEN_1120 = 2'h3 == opidx ? 5'h7 : 5'h0; // @[NulCtrlMP.scala 370:{28,28} 47:30]
  wire [63:0] _GEN_1121 = 2'h0 == opidx ? 64'h1f : 64'h0; // @[NulCtrlMP.scala 371:{30,30} 48:32]
  wire [63:0] _GEN_1122 = 2'h1 == opidx ? 64'h1f : 64'h0; // @[NulCtrlMP.scala 371:{30,30} 48:32]
  wire [63:0] _GEN_1123 = 2'h2 == opidx ? 64'h1f : 64'h0; // @[NulCtrlMP.scala 371:{30,30} 48:32]
  wire [63:0] _GEN_1124 = 2'h3 == opidx ? 64'h1f : 64'h0; // @[NulCtrlMP.scala 371:{30,30} 48:32]
  wire  _GEN_1126 = 2'h1 == opidx ? io_cpu_1_regacc_busy : io_cpu_0_regacc_busy; // @[NulCtrlMP.scala 372:{14,14}]
  wire  _GEN_1127 = 2'h2 == opidx ? io_cpu_2_regacc_busy : _GEN_1126; // @[NulCtrlMP.scala 372:{14,14}]
  wire  _GEN_1128 = 2'h3 == opidx ? io_cpu_3_regacc_busy : _GEN_1127; // @[NulCtrlMP.scala 372:{14,14}]
  wire  _T_122 = ~_GEN_1128; // @[NulCtrlMP.scala 372:14]
  wire [128:0] _GEN_1129 = ~_GEN_1128 ? _cnt_T : _GEN_1112; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_1130 = cnt[1] & _GEN_145; // @[NulCtrlMP.scala 423:22 46:29]
  wire  _GEN_1131 = cnt[1] & _GEN_146; // @[NulCtrlMP.scala 423:22 46:29]
  wire  _GEN_1132 = cnt[1] & _GEN_147; // @[NulCtrlMP.scala 423:22 46:29]
  wire  _GEN_1133 = cnt[1] & _GEN_148; // @[NulCtrlMP.scala 423:22 46:29]
  wire [4:0] _GEN_1134 = cnt[1] ? _GEN_1117 : 5'h0; // @[NulCtrlMP.scala 423:22 47:30]
  wire [4:0] _GEN_1135 = cnt[1] ? _GEN_1118 : 5'h0; // @[NulCtrlMP.scala 423:22 47:30]
  wire [4:0] _GEN_1136 = cnt[1] ? _GEN_1119 : 5'h0; // @[NulCtrlMP.scala 423:22 47:30]
  wire [4:0] _GEN_1137 = cnt[1] ? _GEN_1120 : 5'h0; // @[NulCtrlMP.scala 423:22 47:30]
  wire [63:0] _GEN_1138 = cnt[1] ? _GEN_1121 : 64'h0; // @[NulCtrlMP.scala 423:22 48:32]
  wire [63:0] _GEN_1139 = cnt[1] ? _GEN_1122 : 64'h0; // @[NulCtrlMP.scala 423:22 48:32]
  wire [63:0] _GEN_1140 = cnt[1] ? _GEN_1123 : 64'h0; // @[NulCtrlMP.scala 423:22 48:32]
  wire [63:0] _GEN_1141 = cnt[1] ? _GEN_1124 : 64'h0; // @[NulCtrlMP.scala 423:22 48:32]
  wire [128:0] _GEN_1142 = cnt[1] ? _GEN_1129 : _GEN_1112; // @[NulCtrlMP.scala 423:22]
  wire  _GEN_1143 = _GEN_145 | _GEN_1130; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1144 = _GEN_146 | _GEN_1131; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1145 = _GEN_147 | _GEN_1132; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1146 = _GEN_148 | _GEN_1133; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_1147 = 2'h0 == opidx ? 5'h8 : _GEN_1134; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1148 = 2'h1 == opidx ? 5'h8 : _GEN_1135; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1149 = 2'h2 == opidx ? 5'h8 : _GEN_1136; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1150 = 2'h3 == opidx ? 5'h8 : _GEN_1137; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_1151 = 2'h0 == opidx ? 64'h7fffffffff : _GEN_1138; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1152 = 2'h1 == opidx ? 64'h7fffffffff : _GEN_1139; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1153 = 2'h2 == opidx ? 64'h7fffffffff : _GEN_1140; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1154 = 2'h3 == opidx ? 64'h7fffffffff : _GEN_1141; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_1155 = ~_GEN_1128 ? _cnt_T : _GEN_1142; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_1156 = cnt[2] ? _GEN_1143 : _GEN_1130; // @[NulCtrlMP.scala 424:22]
  wire  _GEN_1157 = cnt[2] ? _GEN_1144 : _GEN_1131; // @[NulCtrlMP.scala 424:22]
  wire  _GEN_1158 = cnt[2] ? _GEN_1145 : _GEN_1132; // @[NulCtrlMP.scala 424:22]
  wire  _GEN_1159 = cnt[2] ? _GEN_1146 : _GEN_1133; // @[NulCtrlMP.scala 424:22]
  wire [4:0] _GEN_1160 = cnt[2] ? _GEN_1147 : _GEN_1134; // @[NulCtrlMP.scala 424:22]
  wire [4:0] _GEN_1161 = cnt[2] ? _GEN_1148 : _GEN_1135; // @[NulCtrlMP.scala 424:22]
  wire [4:0] _GEN_1162 = cnt[2] ? _GEN_1149 : _GEN_1136; // @[NulCtrlMP.scala 424:22]
  wire [4:0] _GEN_1163 = cnt[2] ? _GEN_1150 : _GEN_1137; // @[NulCtrlMP.scala 424:22]
  wire [63:0] _GEN_1164 = cnt[2] ? _GEN_1151 : _GEN_1138; // @[NulCtrlMP.scala 424:22]
  wire [63:0] _GEN_1165 = cnt[2] ? _GEN_1152 : _GEN_1139; // @[NulCtrlMP.scala 424:22]
  wire [63:0] _GEN_1166 = cnt[2] ? _GEN_1153 : _GEN_1140; // @[NulCtrlMP.scala 424:22]
  wire [63:0] _GEN_1167 = cnt[2] ? _GEN_1154 : _GEN_1141; // @[NulCtrlMP.scala 424:22]
  wire [128:0] _GEN_1168 = cnt[2] ? _GEN_1155 : _GEN_1142; // @[NulCtrlMP.scala 424:22]
  wire [31:0] _GEN_1173 = 2'h0 == opidx ? 32'h3a039073 : 32'h0; // @[NulCtrlMP.scala 395:{28,28} 50:30]
  wire [31:0] _GEN_1174 = 2'h1 == opidx ? 32'h3a039073 : 32'h0; // @[NulCtrlMP.scala 395:{28,28} 50:30]
  wire [31:0] _GEN_1175 = 2'h2 == opidx ? 32'h3a039073 : 32'h0; // @[NulCtrlMP.scala 395:{28,28} 50:30]
  wire [31:0] _GEN_1176 = 2'h3 == opidx ? 32'h3a039073 : 32'h0; // @[NulCtrlMP.scala 395:{28,28} 50:30]
  wire  _GEN_1178 = 2'h1 == opidx ? io_cpu_1_inst64_ready : io_cpu_0_inst64_ready; // @[NulCtrlMP.scala 396:{36,36}]
  wire  _GEN_1179 = 2'h2 == opidx ? io_cpu_2_inst64_ready : _GEN_1178; // @[NulCtrlMP.scala 396:{36,36}]
  wire  _GEN_1180 = 2'h3 == opidx ? io_cpu_3_inst64_ready : _GEN_1179; // @[NulCtrlMP.scala 396:{36,36}]
  wire [128:0] _GEN_1181 = _GEN_1180 ? _cnt_T : _GEN_1168; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1182 = cnt[3] & _GEN_145; // @[NulCtrlMP.scala 425:22 49:26]
  wire  _GEN_1183 = cnt[3] & _GEN_146; // @[NulCtrlMP.scala 425:22 49:26]
  wire  _GEN_1184 = cnt[3] & _GEN_147; // @[NulCtrlMP.scala 425:22 49:26]
  wire  _GEN_1185 = cnt[3] & _GEN_148; // @[NulCtrlMP.scala 425:22 49:26]
  wire [31:0] _GEN_1186 = cnt[3] ? _GEN_1173 : 32'h0; // @[NulCtrlMP.scala 425:22 50:30]
  wire [31:0] _GEN_1187 = cnt[3] ? _GEN_1174 : 32'h0; // @[NulCtrlMP.scala 425:22 50:30]
  wire [31:0] _GEN_1188 = cnt[3] ? _GEN_1175 : 32'h0; // @[NulCtrlMP.scala 425:22 50:30]
  wire [31:0] _GEN_1189 = cnt[3] ? _GEN_1176 : 32'h0; // @[NulCtrlMP.scala 425:22 50:30]
  wire [128:0] _GEN_1190 = cnt[3] ? _GEN_1181 : _GEN_1168; // @[NulCtrlMP.scala 425:22]
  wire  _GEN_1191 = _GEN_145 | _GEN_1182; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1192 = _GEN_146 | _GEN_1183; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1193 = _GEN_147 | _GEN_1184; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1194 = _GEN_148 | _GEN_1185; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_1195 = 2'h0 == opidx ? 32'h3b041073 : _GEN_1186; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1196 = 2'h1 == opidx ? 32'h3b041073 : _GEN_1187; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1197 = 2'h2 == opidx ? 32'h3b041073 : _GEN_1188; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1198 = 2'h3 == opidx ? 32'h3b041073 : _GEN_1189; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_1199 = _GEN_1180 ? _cnt_T : _GEN_1190; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1200 = cnt[4] ? _GEN_1191 : _GEN_1182; // @[NulCtrlMP.scala 426:22]
  wire  _GEN_1201 = cnt[4] ? _GEN_1192 : _GEN_1183; // @[NulCtrlMP.scala 426:22]
  wire  _GEN_1202 = cnt[4] ? _GEN_1193 : _GEN_1184; // @[NulCtrlMP.scala 426:22]
  wire  _GEN_1203 = cnt[4] ? _GEN_1194 : _GEN_1185; // @[NulCtrlMP.scala 426:22]
  wire [31:0] _GEN_1204 = cnt[4] ? _GEN_1195 : _GEN_1186; // @[NulCtrlMP.scala 426:22]
  wire [31:0] _GEN_1205 = cnt[4] ? _GEN_1196 : _GEN_1187; // @[NulCtrlMP.scala 426:22]
  wire [31:0] _GEN_1206 = cnt[4] ? _GEN_1197 : _GEN_1188; // @[NulCtrlMP.scala 426:22]
  wire [31:0] _GEN_1207 = cnt[4] ? _GEN_1198 : _GEN_1189; // @[NulCtrlMP.scala 426:22]
  wire [128:0] _GEN_1208 = cnt[4] ? _GEN_1199 : _GEN_1190; // @[NulCtrlMP.scala 426:22]
  wire  _GEN_1209 = _GEN_145 | _GEN_1200; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1210 = _GEN_146 | _GEN_1201; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1211 = _GEN_147 | _GEN_1202; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1212 = _GEN_148 | _GEN_1203; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_1213 = 2'h0 == opidx ? 32'h22b7 : _GEN_1204; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1214 = 2'h1 == opidx ? 32'h22b7 : _GEN_1205; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1215 = 2'h2 == opidx ? 32'h22b7 : _GEN_1206; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1216 = 2'h3 == opidx ? 32'h22b7 : _GEN_1207; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_1217 = _GEN_1180 ? _cnt_T : _GEN_1208; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1218 = cnt[5] ? _GEN_1209 : _GEN_1200; // @[NulCtrlMP.scala 427:22]
  wire  _GEN_1219 = cnt[5] ? _GEN_1210 : _GEN_1201; // @[NulCtrlMP.scala 427:22]
  wire  _GEN_1220 = cnt[5] ? _GEN_1211 : _GEN_1202; // @[NulCtrlMP.scala 427:22]
  wire  _GEN_1221 = cnt[5] ? _GEN_1212 : _GEN_1203; // @[NulCtrlMP.scala 427:22]
  wire [31:0] _GEN_1222 = cnt[5] ? _GEN_1213 : _GEN_1204; // @[NulCtrlMP.scala 427:22]
  wire [31:0] _GEN_1223 = cnt[5] ? _GEN_1214 : _GEN_1205; // @[NulCtrlMP.scala 427:22]
  wire [31:0] _GEN_1224 = cnt[5] ? _GEN_1215 : _GEN_1206; // @[NulCtrlMP.scala 427:22]
  wire [31:0] _GEN_1225 = cnt[5] ? _GEN_1216 : _GEN_1207; // @[NulCtrlMP.scala 427:22]
  wire [128:0] _GEN_1226 = cnt[5] ? _GEN_1217 : _GEN_1208; // @[NulCtrlMP.scala 427:22]
  wire  _GEN_1227 = _GEN_145 | _GEN_1218; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1228 = _GEN_146 | _GEN_1219; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1229 = _GEN_147 | _GEN_1220; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1230 = _GEN_148 | _GEN_1221; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_1231 = 2'h0 == opidx ? 32'h3002a073 : _GEN_1222; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1232 = 2'h1 == opidx ? 32'h3002a073 : _GEN_1223; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1233 = 2'h2 == opidx ? 32'h3002a073 : _GEN_1224; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1234 = 2'h3 == opidx ? 32'h3002a073 : _GEN_1225; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_1235 = _GEN_1180 ? _cnt_T : _GEN_1226; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1236 = cnt[6] ? _GEN_1227 : _GEN_1218; // @[NulCtrlMP.scala 434:22]
  wire  _GEN_1237 = cnt[6] ? _GEN_1228 : _GEN_1219; // @[NulCtrlMP.scala 434:22]
  wire  _GEN_1238 = cnt[6] ? _GEN_1229 : _GEN_1220; // @[NulCtrlMP.scala 434:22]
  wire  _GEN_1239 = cnt[6] ? _GEN_1230 : _GEN_1221; // @[NulCtrlMP.scala 434:22]
  wire [31:0] _GEN_1240 = cnt[6] ? _GEN_1231 : _GEN_1222; // @[NulCtrlMP.scala 434:22]
  wire [31:0] _GEN_1241 = cnt[6] ? _GEN_1232 : _GEN_1223; // @[NulCtrlMP.scala 434:22]
  wire [31:0] _GEN_1242 = cnt[6] ? _GEN_1233 : _GEN_1224; // @[NulCtrlMP.scala 434:22]
  wire [31:0] _GEN_1243 = cnt[6] ? _GEN_1234 : _GEN_1225; // @[NulCtrlMP.scala 434:22]
  wire [128:0] _GEN_1244 = cnt[6] ? _GEN_1235 : _GEN_1226; // @[NulCtrlMP.scala 434:22]
  wire  _GEN_1250 = 2'h1 == opidx ? io_cpu_1_inst64_busy : io_cpu_0_inst64_busy; // @[NulCtrlMP.scala 402:{14,14}]
  wire  _GEN_1251 = 2'h2 == opidx ? io_cpu_2_inst64_busy : _GEN_1250; // @[NulCtrlMP.scala 402:{14,14}]
  wire  _GEN_1252 = 2'h3 == opidx ? io_cpu_3_inst64_busy : _GEN_1251; // @[NulCtrlMP.scala 402:{14,14}]
  wire [128:0] _GEN_1253 = ~_GEN_1252 ? _cnt_T : _GEN_1244; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_1254 = cnt[7] & _GEN_145; // @[NulCtrlMP.scala 441:22 52:32]
  wire  _GEN_1255 = cnt[7] & _GEN_146; // @[NulCtrlMP.scala 441:22 52:32]
  wire  _GEN_1256 = cnt[7] & _GEN_147; // @[NulCtrlMP.scala 441:22 52:32]
  wire  _GEN_1257 = cnt[7] & _GEN_148; // @[NulCtrlMP.scala 441:22 52:32]
  wire [128:0] _GEN_1258 = cnt[7] ? _GEN_1253 : _GEN_1244; // @[NulCtrlMP.scala 441:22]
  wire [1:0] _nextidx_T_1 = init_cnt + 2'h1; // @[NulCtrlMP.scala 447:41]
  wire [7:0] nextidx = {{6'd0}, _nextidx_T_1}; // @[NulCtrlMP.scala 447:51]
  wire [4:0] _GEN_1259 = init_cnt == 2'h3 ? 5'h1f : _GEN_1111; // @[NulCtrlMP.scala 444:47 445:23]
  wire [128:0] _GEN_1262 = cnt[8] ? 129'h1 : _GEN_1258; // @[NulCtrlMP.scala 442:22 443:17]
  wire [4:0] _GEN_1263 = cnt[8] ? _GEN_1259 : _GEN_1111; // @[NulCtrlMP.scala 442:22]
  wire [128:0] _GEN_1266 = state == 5'h1 ? _GEN_1262 : {{1'd0}, cnt}; // @[NulCtrlMP.scala 345:22 421:35]
  wire  _GEN_1267 = state == 5'h1 & _GEN_1156; // @[NulCtrlMP.scala 421:35 46:29]
  wire  _GEN_1268 = state == 5'h1 & _GEN_1157; // @[NulCtrlMP.scala 421:35 46:29]
  wire  _GEN_1269 = state == 5'h1 & _GEN_1158; // @[NulCtrlMP.scala 421:35 46:29]
  wire  _GEN_1270 = state == 5'h1 & _GEN_1159; // @[NulCtrlMP.scala 421:35 46:29]
  wire [4:0] _GEN_1271 = state == 5'h1 ? _GEN_1160 : 5'h0; // @[NulCtrlMP.scala 421:35 47:30]
  wire [4:0] _GEN_1272 = state == 5'h1 ? _GEN_1161 : 5'h0; // @[NulCtrlMP.scala 421:35 47:30]
  wire [4:0] _GEN_1273 = state == 5'h1 ? _GEN_1162 : 5'h0; // @[NulCtrlMP.scala 421:35 47:30]
  wire [4:0] _GEN_1274 = state == 5'h1 ? _GEN_1163 : 5'h0; // @[NulCtrlMP.scala 421:35 47:30]
  wire [63:0] _GEN_1275 = state == 5'h1 ? _GEN_1164 : 64'h0; // @[NulCtrlMP.scala 421:35 48:32]
  wire [63:0] _GEN_1276 = state == 5'h1 ? _GEN_1165 : 64'h0; // @[NulCtrlMP.scala 421:35 48:32]
  wire [63:0] _GEN_1277 = state == 5'h1 ? _GEN_1166 : 64'h0; // @[NulCtrlMP.scala 421:35 48:32]
  wire [63:0] _GEN_1278 = state == 5'h1 ? _GEN_1167 : 64'h0; // @[NulCtrlMP.scala 421:35 48:32]
  wire  _GEN_1279 = state == 5'h1 & _GEN_1236; // @[NulCtrlMP.scala 421:35 49:26]
  wire  _GEN_1280 = state == 5'h1 & _GEN_1237; // @[NulCtrlMP.scala 421:35 49:26]
  wire  _GEN_1281 = state == 5'h1 & _GEN_1238; // @[NulCtrlMP.scala 421:35 49:26]
  wire  _GEN_1282 = state == 5'h1 & _GEN_1239; // @[NulCtrlMP.scala 421:35 49:26]
  wire [31:0] _GEN_1283 = state == 5'h1 ? _GEN_1240 : 32'h0; // @[NulCtrlMP.scala 421:35 50:30]
  wire [31:0] _GEN_1284 = state == 5'h1 ? _GEN_1241 : 32'h0; // @[NulCtrlMP.scala 421:35 50:30]
  wire [31:0] _GEN_1285 = state == 5'h1 ? _GEN_1242 : 32'h0; // @[NulCtrlMP.scala 421:35 50:30]
  wire [31:0] _GEN_1286 = state == 5'h1 ? _GEN_1243 : 32'h0; // @[NulCtrlMP.scala 421:35 50:30]
  wire  _GEN_1287 = state == 5'h1 & _GEN_1254; // @[NulCtrlMP.scala 421:35 52:32]
  wire  _GEN_1288 = state == 5'h1 & _GEN_1255; // @[NulCtrlMP.scala 421:35 52:32]
  wire  _GEN_1289 = state == 5'h1 & _GEN_1256; // @[NulCtrlMP.scala 421:35 52:32]
  wire  _GEN_1290 = state == 5'h1 & _GEN_1257; // @[NulCtrlMP.scala 421:35 52:32]
  wire [4:0] _GEN_1291 = state == 5'h1 ? _GEN_1263 : _GEN_1111; // @[NulCtrlMP.scala 421:35]
  wire [31:0] _T_135 = {oparg_5,oparg_4,oparg_3,oparg_2}; // @[Cat.scala 31:58]
  wire  _GEN_1294 = _GEN_145 | _GEN_1279; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1295 = _GEN_146 | _GEN_1280; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1296 = _GEN_147 | _GEN_1281; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1297 = _GEN_148 | _GEN_1282; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_1298 = 2'h0 == opidx ? _T_135 : _GEN_1283; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1299 = 2'h1 == opidx ? _T_135 : _GEN_1284; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1300 = 2'h2 == opidx ? _T_135 : _GEN_1285; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1301 = 2'h3 == opidx ? _T_135 : _GEN_1286; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_1302 = _GEN_1180 ? _cnt_T : _GEN_1266; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1303 = cnt[0] ? _GEN_1294 : _GEN_1279; // @[NulCtrlMP.scala 455:22]
  wire  _GEN_1304 = cnt[0] ? _GEN_1295 : _GEN_1280; // @[NulCtrlMP.scala 455:22]
  wire  _GEN_1305 = cnt[0] ? _GEN_1296 : _GEN_1281; // @[NulCtrlMP.scala 455:22]
  wire  _GEN_1306 = cnt[0] ? _GEN_1297 : _GEN_1282; // @[NulCtrlMP.scala 455:22]
  wire [31:0] _GEN_1307 = cnt[0] ? _GEN_1298 : _GEN_1283; // @[NulCtrlMP.scala 455:22]
  wire [31:0] _GEN_1308 = cnt[0] ? _GEN_1299 : _GEN_1284; // @[NulCtrlMP.scala 455:22]
  wire [31:0] _GEN_1309 = cnt[0] ? _GEN_1300 : _GEN_1285; // @[NulCtrlMP.scala 455:22]
  wire [31:0] _GEN_1310 = cnt[0] ? _GEN_1301 : _GEN_1286; // @[NulCtrlMP.scala 455:22]
  wire [128:0] _GEN_1311 = cnt[0] ? _GEN_1302 : _GEN_1266; // @[NulCtrlMP.scala 455:22]
  wire  _GEN_1312 = _GEN_145 | _GEN_1287; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1313 = _GEN_146 | _GEN_1288; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1314 = _GEN_147 | _GEN_1289; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1315 = _GEN_148 | _GEN_1290; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_1316 = ~_GEN_1252 ? _cnt_T : _GEN_1311; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_1317 = cnt[1] ? _GEN_1312 : _GEN_1287; // @[NulCtrlMP.scala 456:22]
  wire  _GEN_1318 = cnt[1] ? _GEN_1313 : _GEN_1288; // @[NulCtrlMP.scala 456:22]
  wire  _GEN_1319 = cnt[1] ? _GEN_1314 : _GEN_1289; // @[NulCtrlMP.scala 456:22]
  wire  _GEN_1320 = cnt[1] ? _GEN_1315 : _GEN_1290; // @[NulCtrlMP.scala 456:22]
  wire [128:0] _GEN_1321 = cnt[1] ? _GEN_1316 : _GEN_1311; // @[NulCtrlMP.scala 456:22]
  wire [128:0] _GEN_1322 = cnt[2] ? 129'h1 : _GEN_1321; // @[NulCtrlMP.scala 457:22 458:17]
  wire [4:0] _GEN_1323 = cnt[2] ? 5'h5 : _GEN_1291; // @[NulCtrlMP.scala 457:22 459:19]
  wire  _GEN_1324 = state == 5'h17 ? _GEN_1303 : _GEN_1279; // @[NulCtrlMP.scala 454:32]
  wire  _GEN_1325 = state == 5'h17 ? _GEN_1304 : _GEN_1280; // @[NulCtrlMP.scala 454:32]
  wire  _GEN_1326 = state == 5'h17 ? _GEN_1305 : _GEN_1281; // @[NulCtrlMP.scala 454:32]
  wire  _GEN_1327 = state == 5'h17 ? _GEN_1306 : _GEN_1282; // @[NulCtrlMP.scala 454:32]
  wire [31:0] _GEN_1328 = state == 5'h17 ? _GEN_1307 : _GEN_1283; // @[NulCtrlMP.scala 454:32]
  wire [31:0] _GEN_1329 = state == 5'h17 ? _GEN_1308 : _GEN_1284; // @[NulCtrlMP.scala 454:32]
  wire [31:0] _GEN_1330 = state == 5'h17 ? _GEN_1309 : _GEN_1285; // @[NulCtrlMP.scala 454:32]
  wire [31:0] _GEN_1331 = state == 5'h17 ? _GEN_1310 : _GEN_1286; // @[NulCtrlMP.scala 454:32]
  wire [128:0] _GEN_1332 = state == 5'h17 ? _GEN_1322 : _GEN_1266; // @[NulCtrlMP.scala 454:32]
  wire  _GEN_1333 = state == 5'h17 ? _GEN_1317 : _GEN_1287; // @[NulCtrlMP.scala 454:32]
  wire  _GEN_1334 = state == 5'h17 ? _GEN_1318 : _GEN_1288; // @[NulCtrlMP.scala 454:32]
  wire  _GEN_1335 = state == 5'h17 ? _GEN_1319 : _GEN_1289; // @[NulCtrlMP.scala 454:32]
  wire  _GEN_1336 = state == 5'h17 ? _GEN_1320 : _GEN_1290; // @[NulCtrlMP.scala 454:32]
  wire [4:0] _GEN_1337 = state == 5'h17 ? _GEN_1323 : _GEN_1291; // @[NulCtrlMP.scala 454:32]
  wire [63:0] satp_value = {4'h8,oparg_3,oparg_2,4'h0,oparg_8,oparg_7,oparg_6,oparg_5,oparg_4}; // @[Cat.scala 31:58]
  wire [4:0] _GEN_1342 = 2'h0 == opidx ? 5'h5 : _GEN_1271; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1343 = 2'h1 == opidx ? 5'h5 : _GEN_1272; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1344 = 2'h2 == opidx ? 5'h5 : _GEN_1273; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1345 = 2'h3 == opidx ? 5'h5 : _GEN_1274; // @[NulCtrlMP.scala 352:{28,28}]
  wire [63:0] _GEN_1347 = 2'h1 == opidx ? io_cpu_1_regacc_rdata : io_cpu_0_regacc_rdata; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_1348 = 2'h2 == opidx ? io_cpu_2_regacc_rdata : _GEN_1347; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_1349 = 2'h3 == opidx ? io_cpu_3_regacc_rdata : _GEN_1348; // @[NulCtrlMP.scala 355:{17,17}]
  wire [128:0] _GEN_1350 = _T_122 ? _cnt_T : _GEN_1332; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_1351 = _T_122 ? _GEN_1349 : regback_0; // @[NulCtrlMP.scala 353:36 355:17 346:26]
  wire  _GEN_1352 = cnt[0] & _GEN_145; // @[NulCtrlMP.scala 408:32 45:29]
  wire  _GEN_1353 = cnt[0] & _GEN_146; // @[NulCtrlMP.scala 408:32 45:29]
  wire  _GEN_1354 = cnt[0] & _GEN_147; // @[NulCtrlMP.scala 408:32 45:29]
  wire  _GEN_1355 = cnt[0] & _GEN_148; // @[NulCtrlMP.scala 408:32 45:29]
  wire [4:0] _GEN_1356 = cnt[0] ? _GEN_1342 : _GEN_1271; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1357 = cnt[0] ? _GEN_1343 : _GEN_1272; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1358 = cnt[0] ? _GEN_1344 : _GEN_1273; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1359 = cnt[0] ? _GEN_1345 : _GEN_1274; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_1360 = cnt[0] ? _GEN_1350 : _GEN_1332; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_1361 = cnt[0] ? _GEN_1351 : regback_0; // @[NulCtrlMP.scala 346:26 408:32]
  wire  _GEN_1362 = _GEN_145 | _GEN_1267; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1363 = _GEN_146 | _GEN_1268; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1364 = _GEN_147 | _GEN_1269; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1365 = _GEN_148 | _GEN_1270; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_1366 = 2'h0 == opidx ? 5'h5 : _GEN_1356; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1367 = 2'h1 == opidx ? 5'h5 : _GEN_1357; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1368 = 2'h2 == opidx ? 5'h5 : _GEN_1358; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1369 = 2'h3 == opidx ? 5'h5 : _GEN_1359; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_1370 = 2'h0 == opidx ? satp_value : _GEN_1275; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1371 = 2'h1 == opidx ? satp_value : _GEN_1276; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1372 = 2'h2 == opidx ? satp_value : _GEN_1277; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1373 = 2'h3 == opidx ? satp_value : _GEN_1278; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_1374 = ~_GEN_1128 ? _cnt_T : _GEN_1360; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_1375 = cnt[1] ? _GEN_1362 : _GEN_1267; // @[NulCtrlMP.scala 478:22]
  wire  _GEN_1376 = cnt[1] ? _GEN_1363 : _GEN_1268; // @[NulCtrlMP.scala 478:22]
  wire  _GEN_1377 = cnt[1] ? _GEN_1364 : _GEN_1269; // @[NulCtrlMP.scala 478:22]
  wire  _GEN_1378 = cnt[1] ? _GEN_1365 : _GEN_1270; // @[NulCtrlMP.scala 478:22]
  wire [4:0] _GEN_1379 = cnt[1] ? _GEN_1366 : _GEN_1356; // @[NulCtrlMP.scala 478:22]
  wire [4:0] _GEN_1380 = cnt[1] ? _GEN_1367 : _GEN_1357; // @[NulCtrlMP.scala 478:22]
  wire [4:0] _GEN_1381 = cnt[1] ? _GEN_1368 : _GEN_1358; // @[NulCtrlMP.scala 478:22]
  wire [4:0] _GEN_1382 = cnt[1] ? _GEN_1369 : _GEN_1359; // @[NulCtrlMP.scala 478:22]
  wire [63:0] _GEN_1383 = cnt[1] ? _GEN_1370 : _GEN_1275; // @[NulCtrlMP.scala 478:22]
  wire [63:0] _GEN_1384 = cnt[1] ? _GEN_1371 : _GEN_1276; // @[NulCtrlMP.scala 478:22]
  wire [63:0] _GEN_1385 = cnt[1] ? _GEN_1372 : _GEN_1277; // @[NulCtrlMP.scala 478:22]
  wire [63:0] _GEN_1386 = cnt[1] ? _GEN_1373 : _GEN_1278; // @[NulCtrlMP.scala 478:22]
  wire [128:0] _GEN_1387 = cnt[1] ? _GEN_1374 : _GEN_1360; // @[NulCtrlMP.scala 478:22]
  wire  _GEN_1388 = _GEN_145 | _GEN_1324; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1389 = _GEN_146 | _GEN_1325; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1390 = _GEN_147 | _GEN_1326; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1391 = _GEN_148 | _GEN_1327; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_1392 = 2'h0 == opidx ? 32'h18029073 : _GEN_1328; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1393 = 2'h1 == opidx ? 32'h18029073 : _GEN_1329; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1394 = 2'h2 == opidx ? 32'h18029073 : _GEN_1330; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1395 = 2'h3 == opidx ? 32'h18029073 : _GEN_1331; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_1396 = _GEN_1180 ? _cnt_T : _GEN_1387; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1397 = cnt[2] ? _GEN_1388 : _GEN_1324; // @[NulCtrlMP.scala 479:22]
  wire  _GEN_1398 = cnt[2] ? _GEN_1389 : _GEN_1325; // @[NulCtrlMP.scala 479:22]
  wire  _GEN_1399 = cnt[2] ? _GEN_1390 : _GEN_1326; // @[NulCtrlMP.scala 479:22]
  wire  _GEN_1400 = cnt[2] ? _GEN_1391 : _GEN_1327; // @[NulCtrlMP.scala 479:22]
  wire [31:0] _GEN_1401 = cnt[2] ? _GEN_1392 : _GEN_1328; // @[NulCtrlMP.scala 479:22]
  wire [31:0] _GEN_1402 = cnt[2] ? _GEN_1393 : _GEN_1329; // @[NulCtrlMP.scala 479:22]
  wire [31:0] _GEN_1403 = cnt[2] ? _GEN_1394 : _GEN_1330; // @[NulCtrlMP.scala 479:22]
  wire [31:0] _GEN_1404 = cnt[2] ? _GEN_1395 : _GEN_1331; // @[NulCtrlMP.scala 479:22]
  wire [128:0] _GEN_1405 = cnt[2] ? _GEN_1396 : _GEN_1387; // @[NulCtrlMP.scala 479:22]
  wire  _GEN_1406 = _GEN_145 | _GEN_1333; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1407 = _GEN_146 | _GEN_1334; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1408 = _GEN_147 | _GEN_1335; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1409 = _GEN_148 | _GEN_1336; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_1410 = ~_GEN_1252 ? _cnt_T : _GEN_1405; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_1411 = cnt[3] ? _GEN_1406 : _GEN_1333; // @[NulCtrlMP.scala 480:22]
  wire  _GEN_1412 = cnt[3] ? _GEN_1407 : _GEN_1334; // @[NulCtrlMP.scala 480:22]
  wire  _GEN_1413 = cnt[3] ? _GEN_1408 : _GEN_1335; // @[NulCtrlMP.scala 480:22]
  wire  _GEN_1414 = cnt[3] ? _GEN_1409 : _GEN_1336; // @[NulCtrlMP.scala 480:22]
  wire [128:0] _GEN_1415 = cnt[3] ? _GEN_1410 : _GEN_1405; // @[NulCtrlMP.scala 480:22]
  wire  _GEN_1416 = _GEN_145 | _GEN_1375; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1417 = _GEN_146 | _GEN_1376; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1418 = _GEN_147 | _GEN_1377; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1419 = _GEN_148 | _GEN_1378; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_1420 = 2'h0 == opidx ? 5'h5 : _GEN_1379; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1421 = 2'h1 == opidx ? 5'h5 : _GEN_1380; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1422 = 2'h2 == opidx ? 5'h5 : _GEN_1381; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1423 = 2'h3 == opidx ? 5'h5 : _GEN_1382; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_1424 = 2'h0 == opidx ? regback_0 : _GEN_1383; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1425 = 2'h1 == opidx ? regback_0 : _GEN_1384; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1426 = 2'h2 == opidx ? regback_0 : _GEN_1385; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1427 = 2'h3 == opidx ? regback_0 : _GEN_1386; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_1428 = ~_GEN_1128 ? _cnt_T : _GEN_1415; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_1429 = cnt[4] ? _GEN_1416 : _GEN_1375; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1430 = cnt[4] ? _GEN_1417 : _GEN_1376; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1431 = cnt[4] ? _GEN_1418 : _GEN_1377; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1432 = cnt[4] ? _GEN_1419 : _GEN_1378; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1433 = cnt[4] ? _GEN_1420 : _GEN_1379; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1434 = cnt[4] ? _GEN_1421 : _GEN_1380; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1435 = cnt[4] ? _GEN_1422 : _GEN_1381; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1436 = cnt[4] ? _GEN_1423 : _GEN_1382; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1437 = cnt[4] ? _GEN_1424 : _GEN_1383; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1438 = cnt[4] ? _GEN_1425 : _GEN_1384; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1439 = cnt[4] ? _GEN_1426 : _GEN_1385; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1440 = cnt[4] ? _GEN_1427 : _GEN_1386; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_1441 = cnt[4] ? _GEN_1428 : _GEN_1415; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_1442 = cnt[5] ? 129'h1 : _GEN_1441; // @[NulCtrlMP.scala 482:22 483:17]
  wire [4:0] _GEN_1443 = cnt[5] ? 5'h5 : _GEN_1337; // @[NulCtrlMP.scala 482:22 484:19]
  wire  _GEN_1444 = state == 5'ha & _GEN_1352; // @[NulCtrlMP.scala 45:29 476:31]
  wire  _GEN_1445 = state == 5'ha & _GEN_1353; // @[NulCtrlMP.scala 45:29 476:31]
  wire  _GEN_1446 = state == 5'ha & _GEN_1354; // @[NulCtrlMP.scala 45:29 476:31]
  wire  _GEN_1447 = state == 5'ha & _GEN_1355; // @[NulCtrlMP.scala 45:29 476:31]
  wire [4:0] _GEN_1448 = state == 5'ha ? _GEN_1433 : _GEN_1271; // @[NulCtrlMP.scala 476:31]
  wire [4:0] _GEN_1449 = state == 5'ha ? _GEN_1434 : _GEN_1272; // @[NulCtrlMP.scala 476:31]
  wire [4:0] _GEN_1450 = state == 5'ha ? _GEN_1435 : _GEN_1273; // @[NulCtrlMP.scala 476:31]
  wire [4:0] _GEN_1451 = state == 5'ha ? _GEN_1436 : _GEN_1274; // @[NulCtrlMP.scala 476:31]
  wire [128:0] _GEN_1452 = state == 5'ha ? _GEN_1442 : _GEN_1332; // @[NulCtrlMP.scala 476:31]
  wire [63:0] _GEN_1453 = state == 5'ha ? _GEN_1361 : regback_0; // @[NulCtrlMP.scala 346:26 476:31]
  wire  _GEN_1454 = state == 5'ha ? _GEN_1429 : _GEN_1267; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1455 = state == 5'ha ? _GEN_1430 : _GEN_1268; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1456 = state == 5'ha ? _GEN_1431 : _GEN_1269; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1457 = state == 5'ha ? _GEN_1432 : _GEN_1270; // @[NulCtrlMP.scala 476:31]
  wire [63:0] _GEN_1458 = state == 5'ha ? _GEN_1437 : _GEN_1275; // @[NulCtrlMP.scala 476:31]
  wire [63:0] _GEN_1459 = state == 5'ha ? _GEN_1438 : _GEN_1276; // @[NulCtrlMP.scala 476:31]
  wire [63:0] _GEN_1460 = state == 5'ha ? _GEN_1439 : _GEN_1277; // @[NulCtrlMP.scala 476:31]
  wire [63:0] _GEN_1461 = state == 5'ha ? _GEN_1440 : _GEN_1278; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1462 = state == 5'ha ? _GEN_1397 : _GEN_1324; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1463 = state == 5'ha ? _GEN_1398 : _GEN_1325; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1464 = state == 5'ha ? _GEN_1399 : _GEN_1326; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1465 = state == 5'ha ? _GEN_1400 : _GEN_1327; // @[NulCtrlMP.scala 476:31]
  wire [31:0] _GEN_1466 = state == 5'ha ? _GEN_1401 : _GEN_1328; // @[NulCtrlMP.scala 476:31]
  wire [31:0] _GEN_1467 = state == 5'ha ? _GEN_1402 : _GEN_1329; // @[NulCtrlMP.scala 476:31]
  wire [31:0] _GEN_1468 = state == 5'ha ? _GEN_1403 : _GEN_1330; // @[NulCtrlMP.scala 476:31]
  wire [31:0] _GEN_1469 = state == 5'ha ? _GEN_1404 : _GEN_1331; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1470 = state == 5'ha ? _GEN_1411 : _GEN_1333; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1471 = state == 5'ha ? _GEN_1412 : _GEN_1334; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1472 = state == 5'ha ? _GEN_1413 : _GEN_1335; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1473 = state == 5'ha ? _GEN_1414 : _GEN_1336; // @[NulCtrlMP.scala 476:31]
  wire [4:0] _GEN_1474 = state == 5'ha ? _GEN_1443 : _GEN_1337; // @[NulCtrlMP.scala 476:31]
  wire  _GEN_1475 = _GEN_145 | _GEN_1462; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1476 = _GEN_146 | _GEN_1463; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1477 = _GEN_147 | _GEN_1464; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1478 = _GEN_148 | _GEN_1465; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_1479 = 2'h0 == opidx ? 32'h12000073 : _GEN_1466; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1480 = 2'h1 == opidx ? 32'h12000073 : _GEN_1467; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1481 = 2'h2 == opidx ? 32'h12000073 : _GEN_1468; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1482 = 2'h3 == opidx ? 32'h12000073 : _GEN_1469; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_1483 = _GEN_1180 ? _cnt_T : _GEN_1452; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1484 = cnt[0] ? _GEN_1475 : _GEN_1462; // @[NulCtrlMP.scala 489:22]
  wire  _GEN_1485 = cnt[0] ? _GEN_1476 : _GEN_1463; // @[NulCtrlMP.scala 489:22]
  wire  _GEN_1486 = cnt[0] ? _GEN_1477 : _GEN_1464; // @[NulCtrlMP.scala 489:22]
  wire  _GEN_1487 = cnt[0] ? _GEN_1478 : _GEN_1465; // @[NulCtrlMP.scala 489:22]
  wire [31:0] _GEN_1488 = cnt[0] ? _GEN_1479 : _GEN_1466; // @[NulCtrlMP.scala 489:22]
  wire [31:0] _GEN_1489 = cnt[0] ? _GEN_1480 : _GEN_1467; // @[NulCtrlMP.scala 489:22]
  wire [31:0] _GEN_1490 = cnt[0] ? _GEN_1481 : _GEN_1468; // @[NulCtrlMP.scala 489:22]
  wire [31:0] _GEN_1491 = cnt[0] ? _GEN_1482 : _GEN_1469; // @[NulCtrlMP.scala 489:22]
  wire [128:0] _GEN_1492 = cnt[0] ? _GEN_1483 : _GEN_1452; // @[NulCtrlMP.scala 489:22]
  wire  _GEN_1493 = _GEN_145 | _GEN_1470; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1494 = _GEN_146 | _GEN_1471; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1495 = _GEN_147 | _GEN_1472; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1496 = _GEN_148 | _GEN_1473; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_1497 = ~_GEN_1252 ? _cnt_T : _GEN_1492; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_1498 = cnt[1] ? _GEN_1493 : _GEN_1470; // @[NulCtrlMP.scala 490:22]
  wire  _GEN_1499 = cnt[1] ? _GEN_1494 : _GEN_1471; // @[NulCtrlMP.scala 490:22]
  wire  _GEN_1500 = cnt[1] ? _GEN_1495 : _GEN_1472; // @[NulCtrlMP.scala 490:22]
  wire  _GEN_1501 = cnt[1] ? _GEN_1496 : _GEN_1473; // @[NulCtrlMP.scala 490:22]
  wire [128:0] _GEN_1502 = cnt[1] ? _GEN_1497 : _GEN_1492; // @[NulCtrlMP.scala 490:22]
  wire [128:0] _GEN_1503 = cnt[2] ? 129'h1 : _GEN_1502; // @[NulCtrlMP.scala 491:22 492:17]
  wire [4:0] _GEN_1504 = cnt[2] ? 5'h5 : _GEN_1474; // @[NulCtrlMP.scala 491:22 493:19]
  wire  _GEN_1505 = state == 5'hc ? _GEN_1484 : _GEN_1462; // @[NulCtrlMP.scala 488:33]
  wire  _GEN_1506 = state == 5'hc ? _GEN_1485 : _GEN_1463; // @[NulCtrlMP.scala 488:33]
  wire  _GEN_1507 = state == 5'hc ? _GEN_1486 : _GEN_1464; // @[NulCtrlMP.scala 488:33]
  wire  _GEN_1508 = state == 5'hc ? _GEN_1487 : _GEN_1465; // @[NulCtrlMP.scala 488:33]
  wire [31:0] _GEN_1509 = state == 5'hc ? _GEN_1488 : _GEN_1466; // @[NulCtrlMP.scala 488:33]
  wire [31:0] _GEN_1510 = state == 5'hc ? _GEN_1489 : _GEN_1467; // @[NulCtrlMP.scala 488:33]
  wire [31:0] _GEN_1511 = state == 5'hc ? _GEN_1490 : _GEN_1468; // @[NulCtrlMP.scala 488:33]
  wire [31:0] _GEN_1512 = state == 5'hc ? _GEN_1491 : _GEN_1469; // @[NulCtrlMP.scala 488:33]
  wire [128:0] _GEN_1513 = state == 5'hc ? _GEN_1503 : _GEN_1452; // @[NulCtrlMP.scala 488:33]
  wire  _GEN_1514 = state == 5'hc ? _GEN_1498 : _GEN_1470; // @[NulCtrlMP.scala 488:33]
  wire  _GEN_1515 = state == 5'hc ? _GEN_1499 : _GEN_1471; // @[NulCtrlMP.scala 488:33]
  wire  _GEN_1516 = state == 5'hc ? _GEN_1500 : _GEN_1472; // @[NulCtrlMP.scala 488:33]
  wire  _GEN_1517 = state == 5'hc ? _GEN_1501 : _GEN_1473; // @[NulCtrlMP.scala 488:33]
  wire [4:0] _GEN_1518 = state == 5'hc ? _GEN_1504 : _GEN_1474; // @[NulCtrlMP.scala 488:33]
  wire [63:0] flush_tlb_address = {12'h0,oparg_8,oparg_7,oparg_6,oparg_5,oparg_4,12'h0}; // @[Cat.scala 31:58]
  wire [16:0] flush_asid = {1'h0,oparg_3,oparg_2}; // @[Cat.scala 31:58]
  wire  _GEN_1519 = _GEN_145 | _GEN_1444; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1520 = _GEN_146 | _GEN_1445; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1521 = _GEN_147 | _GEN_1446; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1522 = _GEN_148 | _GEN_1447; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_1523 = 2'h0 == opidx ? 5'h5 : _GEN_1448; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1524 = 2'h1 == opidx ? 5'h5 : _GEN_1449; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1525 = 2'h2 == opidx ? 5'h5 : _GEN_1450; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1526 = 2'h3 == opidx ? 5'h5 : _GEN_1451; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_1527 = _T_122 ? _cnt_T : _GEN_1513; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_1528 = _T_122 ? _GEN_1349 : _GEN_1453; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_1529 = cnt[0] ? _GEN_1519 : _GEN_1444; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1530 = cnt[0] ? _GEN_1520 : _GEN_1445; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1531 = cnt[0] ? _GEN_1521 : _GEN_1446; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1532 = cnt[0] ? _GEN_1522 : _GEN_1447; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1533 = cnt[0] ? _GEN_1523 : _GEN_1448; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1534 = cnt[0] ? _GEN_1524 : _GEN_1449; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1535 = cnt[0] ? _GEN_1525 : _GEN_1450; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1536 = cnt[0] ? _GEN_1526 : _GEN_1451; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_1537 = cnt[0] ? _GEN_1527 : _GEN_1513; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_1538 = cnt[0] ? _GEN_1528 : _GEN_1453; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1539 = _GEN_145 | _GEN_1529; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1540 = _GEN_146 | _GEN_1530; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1541 = _GEN_147 | _GEN_1531; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1542 = _GEN_148 | _GEN_1532; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_1543 = 2'h0 == opidx ? 5'h6 : _GEN_1533; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1544 = 2'h1 == opidx ? 5'h6 : _GEN_1534; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1545 = 2'h2 == opidx ? 5'h6 : _GEN_1535; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1546 = 2'h3 == opidx ? 5'h6 : _GEN_1536; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_1547 = _T_122 ? _cnt_T : _GEN_1537; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_1548 = _T_122 ? _GEN_1349 : regback_1; // @[NulCtrlMP.scala 353:36 355:17 346:26]
  wire  _GEN_1549 = cnt[1] ? _GEN_1539 : _GEN_1529; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1550 = cnt[1] ? _GEN_1540 : _GEN_1530; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1551 = cnt[1] ? _GEN_1541 : _GEN_1531; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1552 = cnt[1] ? _GEN_1542 : _GEN_1532; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1553 = cnt[1] ? _GEN_1543 : _GEN_1533; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1554 = cnt[1] ? _GEN_1544 : _GEN_1534; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1555 = cnt[1] ? _GEN_1545 : _GEN_1535; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1556 = cnt[1] ? _GEN_1546 : _GEN_1536; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_1557 = cnt[1] ? _GEN_1547 : _GEN_1537; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_1558 = cnt[1] ? _GEN_1548 : regback_1; // @[NulCtrlMP.scala 346:26 408:32]
  wire  _GEN_1559 = _GEN_145 | _GEN_1454; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1560 = _GEN_146 | _GEN_1455; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1561 = _GEN_147 | _GEN_1456; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1562 = _GEN_148 | _GEN_1457; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_1563 = 2'h0 == opidx ? 5'h5 : _GEN_1553; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1564 = 2'h1 == opidx ? 5'h5 : _GEN_1554; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1565 = 2'h2 == opidx ? 5'h5 : _GEN_1555; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1566 = 2'h3 == opidx ? 5'h5 : _GEN_1556; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_1567 = 2'h0 == opidx ? flush_tlb_address : _GEN_1458; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1568 = 2'h1 == opidx ? flush_tlb_address : _GEN_1459; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1569 = 2'h2 == opidx ? flush_tlb_address : _GEN_1460; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1570 = 2'h3 == opidx ? flush_tlb_address : _GEN_1461; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_1571 = ~_GEN_1128 ? _cnt_T : _GEN_1557; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_1572 = cnt[2] ? _GEN_1559 : _GEN_1454; // @[NulCtrlMP.scala 501:22]
  wire  _GEN_1573 = cnt[2] ? _GEN_1560 : _GEN_1455; // @[NulCtrlMP.scala 501:22]
  wire  _GEN_1574 = cnt[2] ? _GEN_1561 : _GEN_1456; // @[NulCtrlMP.scala 501:22]
  wire  _GEN_1575 = cnt[2] ? _GEN_1562 : _GEN_1457; // @[NulCtrlMP.scala 501:22]
  wire [4:0] _GEN_1576 = cnt[2] ? _GEN_1563 : _GEN_1553; // @[NulCtrlMP.scala 501:22]
  wire [4:0] _GEN_1577 = cnt[2] ? _GEN_1564 : _GEN_1554; // @[NulCtrlMP.scala 501:22]
  wire [4:0] _GEN_1578 = cnt[2] ? _GEN_1565 : _GEN_1555; // @[NulCtrlMP.scala 501:22]
  wire [4:0] _GEN_1579 = cnt[2] ? _GEN_1566 : _GEN_1556; // @[NulCtrlMP.scala 501:22]
  wire [63:0] _GEN_1580 = cnt[2] ? _GEN_1567 : _GEN_1458; // @[NulCtrlMP.scala 501:22]
  wire [63:0] _GEN_1581 = cnt[2] ? _GEN_1568 : _GEN_1459; // @[NulCtrlMP.scala 501:22]
  wire [63:0] _GEN_1582 = cnt[2] ? _GEN_1569 : _GEN_1460; // @[NulCtrlMP.scala 501:22]
  wire [63:0] _GEN_1583 = cnt[2] ? _GEN_1570 : _GEN_1461; // @[NulCtrlMP.scala 501:22]
  wire [128:0] _GEN_1584 = cnt[2] ? _GEN_1571 : _GEN_1557; // @[NulCtrlMP.scala 501:22]
  wire  _GEN_1585 = _GEN_145 | _GEN_1572; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1586 = _GEN_146 | _GEN_1573; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1587 = _GEN_147 | _GEN_1574; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1588 = _GEN_148 | _GEN_1575; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_1589 = 2'h0 == opidx ? 5'h6 : _GEN_1576; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1590 = 2'h1 == opidx ? 5'h6 : _GEN_1577; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1591 = 2'h2 == opidx ? 5'h6 : _GEN_1578; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1592 = 2'h3 == opidx ? 5'h6 : _GEN_1579; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _io_cpu_opidx_regacc_wdata_4 = {{47'd0}, flush_asid}; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1593 = 2'h0 == opidx ? _io_cpu_opidx_regacc_wdata_4 : _GEN_1580; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1594 = 2'h1 == opidx ? _io_cpu_opidx_regacc_wdata_4 : _GEN_1581; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1595 = 2'h2 == opidx ? _io_cpu_opidx_regacc_wdata_4 : _GEN_1582; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1596 = 2'h3 == opidx ? _io_cpu_opidx_regacc_wdata_4 : _GEN_1583; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_1597 = ~_GEN_1128 ? _cnt_T : _GEN_1584; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_1598 = cnt[3] ? _GEN_1585 : _GEN_1572; // @[NulCtrlMP.scala 502:22]
  wire  _GEN_1599 = cnt[3] ? _GEN_1586 : _GEN_1573; // @[NulCtrlMP.scala 502:22]
  wire  _GEN_1600 = cnt[3] ? _GEN_1587 : _GEN_1574; // @[NulCtrlMP.scala 502:22]
  wire  _GEN_1601 = cnt[3] ? _GEN_1588 : _GEN_1575; // @[NulCtrlMP.scala 502:22]
  wire [4:0] _GEN_1602 = cnt[3] ? _GEN_1589 : _GEN_1576; // @[NulCtrlMP.scala 502:22]
  wire [4:0] _GEN_1603 = cnt[3] ? _GEN_1590 : _GEN_1577; // @[NulCtrlMP.scala 502:22]
  wire [4:0] _GEN_1604 = cnt[3] ? _GEN_1591 : _GEN_1578; // @[NulCtrlMP.scala 502:22]
  wire [4:0] _GEN_1605 = cnt[3] ? _GEN_1592 : _GEN_1579; // @[NulCtrlMP.scala 502:22]
  wire [63:0] _GEN_1606 = cnt[3] ? _GEN_1593 : _GEN_1580; // @[NulCtrlMP.scala 502:22]
  wire [63:0] _GEN_1607 = cnt[3] ? _GEN_1594 : _GEN_1581; // @[NulCtrlMP.scala 502:22]
  wire [63:0] _GEN_1608 = cnt[3] ? _GEN_1595 : _GEN_1582; // @[NulCtrlMP.scala 502:22]
  wire [63:0] _GEN_1609 = cnt[3] ? _GEN_1596 : _GEN_1583; // @[NulCtrlMP.scala 502:22]
  wire [128:0] _GEN_1610 = cnt[3] ? _GEN_1597 : _GEN_1584; // @[NulCtrlMP.scala 502:22]
  wire  _GEN_1611 = _GEN_145 | _GEN_1505; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1612 = _GEN_146 | _GEN_1506; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1613 = _GEN_147 | _GEN_1507; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1614 = _GEN_148 | _GEN_1508; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_1615 = 2'h0 == opidx ? 32'h12628073 : _GEN_1509; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1616 = 2'h1 == opidx ? 32'h12628073 : _GEN_1510; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1617 = 2'h2 == opidx ? 32'h12628073 : _GEN_1511; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1618 = 2'h3 == opidx ? 32'h12628073 : _GEN_1512; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_1619 = _GEN_1180 ? _cnt_T : _GEN_1610; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1620 = cnt[4] ? _GEN_1611 : _GEN_1505; // @[NulCtrlMP.scala 503:22]
  wire  _GEN_1621 = cnt[4] ? _GEN_1612 : _GEN_1506; // @[NulCtrlMP.scala 503:22]
  wire  _GEN_1622 = cnt[4] ? _GEN_1613 : _GEN_1507; // @[NulCtrlMP.scala 503:22]
  wire  _GEN_1623 = cnt[4] ? _GEN_1614 : _GEN_1508; // @[NulCtrlMP.scala 503:22]
  wire [31:0] _GEN_1624 = cnt[4] ? _GEN_1615 : _GEN_1509; // @[NulCtrlMP.scala 503:22]
  wire [31:0] _GEN_1625 = cnt[4] ? _GEN_1616 : _GEN_1510; // @[NulCtrlMP.scala 503:22]
  wire [31:0] _GEN_1626 = cnt[4] ? _GEN_1617 : _GEN_1511; // @[NulCtrlMP.scala 503:22]
  wire [31:0] _GEN_1627 = cnt[4] ? _GEN_1618 : _GEN_1512; // @[NulCtrlMP.scala 503:22]
  wire [128:0] _GEN_1628 = cnt[4] ? _GEN_1619 : _GEN_1610; // @[NulCtrlMP.scala 503:22]
  wire  _GEN_1629 = _GEN_145 | _GEN_1514; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1630 = _GEN_146 | _GEN_1515; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1631 = _GEN_147 | _GEN_1516; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1632 = _GEN_148 | _GEN_1517; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_1633 = ~_GEN_1252 ? _cnt_T : _GEN_1628; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_1634 = cnt[5] ? _GEN_1629 : _GEN_1514; // @[NulCtrlMP.scala 504:22]
  wire  _GEN_1635 = cnt[5] ? _GEN_1630 : _GEN_1515; // @[NulCtrlMP.scala 504:22]
  wire  _GEN_1636 = cnt[5] ? _GEN_1631 : _GEN_1516; // @[NulCtrlMP.scala 504:22]
  wire  _GEN_1637 = cnt[5] ? _GEN_1632 : _GEN_1517; // @[NulCtrlMP.scala 504:22]
  wire [128:0] _GEN_1638 = cnt[5] ? _GEN_1633 : _GEN_1628; // @[NulCtrlMP.scala 504:22]
  wire  _GEN_1639 = _GEN_145 | _GEN_1598; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1640 = _GEN_146 | _GEN_1599; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1641 = _GEN_147 | _GEN_1600; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1642 = _GEN_148 | _GEN_1601; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_1643 = 2'h0 == opidx ? 5'h5 : _GEN_1602; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1644 = 2'h1 == opidx ? 5'h5 : _GEN_1603; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1645 = 2'h2 == opidx ? 5'h5 : _GEN_1604; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1646 = 2'h3 == opidx ? 5'h5 : _GEN_1605; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_1647 = 2'h0 == opidx ? regback_0 : _GEN_1606; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1648 = 2'h1 == opidx ? regback_0 : _GEN_1607; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1649 = 2'h2 == opidx ? regback_0 : _GEN_1608; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1650 = 2'h3 == opidx ? regback_0 : _GEN_1609; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_1651 = ~_GEN_1128 ? _cnt_T : _GEN_1638; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_1652 = cnt[6] ? _GEN_1639 : _GEN_1598; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1653 = cnt[6] ? _GEN_1640 : _GEN_1599; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1654 = cnt[6] ? _GEN_1641 : _GEN_1600; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1655 = cnt[6] ? _GEN_1642 : _GEN_1601; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1656 = cnt[6] ? _GEN_1643 : _GEN_1602; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1657 = cnt[6] ? _GEN_1644 : _GEN_1603; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1658 = cnt[6] ? _GEN_1645 : _GEN_1604; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1659 = cnt[6] ? _GEN_1646 : _GEN_1605; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1660 = cnt[6] ? _GEN_1647 : _GEN_1606; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1661 = cnt[6] ? _GEN_1648 : _GEN_1607; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1662 = cnt[6] ? _GEN_1649 : _GEN_1608; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1663 = cnt[6] ? _GEN_1650 : _GEN_1609; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_1664 = cnt[6] ? _GEN_1651 : _GEN_1638; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1665 = _GEN_145 | _GEN_1652; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1666 = _GEN_146 | _GEN_1653; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1667 = _GEN_147 | _GEN_1654; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1668 = _GEN_148 | _GEN_1655; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_1669 = 2'h0 == opidx ? 5'h6 : _GEN_1656; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1670 = 2'h1 == opidx ? 5'h6 : _GEN_1657; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1671 = 2'h2 == opidx ? 5'h6 : _GEN_1658; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1672 = 2'h3 == opidx ? 5'h6 : _GEN_1659; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_1673 = 2'h0 == opidx ? regback_1 : _GEN_1660; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1674 = 2'h1 == opidx ? regback_1 : _GEN_1661; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1675 = 2'h2 == opidx ? regback_1 : _GEN_1662; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1676 = 2'h3 == opidx ? regback_1 : _GEN_1663; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_1677 = ~_GEN_1128 ? _cnt_T : _GEN_1664; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_1678 = cnt[7] ? _GEN_1665 : _GEN_1652; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1679 = cnt[7] ? _GEN_1666 : _GEN_1653; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1680 = cnt[7] ? _GEN_1667 : _GEN_1654; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1681 = cnt[7] ? _GEN_1668 : _GEN_1655; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1682 = cnt[7] ? _GEN_1669 : _GEN_1656; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1683 = cnt[7] ? _GEN_1670 : _GEN_1657; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1684 = cnt[7] ? _GEN_1671 : _GEN_1658; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1685 = cnt[7] ? _GEN_1672 : _GEN_1659; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1686 = cnt[7] ? _GEN_1673 : _GEN_1660; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1687 = cnt[7] ? _GEN_1674 : _GEN_1661; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1688 = cnt[7] ? _GEN_1675 : _GEN_1662; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1689 = cnt[7] ? _GEN_1676 : _GEN_1663; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_1690 = cnt[7] ? _GEN_1677 : _GEN_1664; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_1691 = cnt[8] ? 129'h1 : _GEN_1690; // @[NulCtrlMP.scala 506:22 507:17]
  wire [4:0] _GEN_1692 = cnt[8] ? 5'h5 : _GEN_1518; // @[NulCtrlMP.scala 506:22 508:19]
  wire  _GEN_1693 = state == 5'hd ? _GEN_1549 : _GEN_1444; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1694 = state == 5'hd ? _GEN_1550 : _GEN_1445; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1695 = state == 5'hd ? _GEN_1551 : _GEN_1446; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1696 = state == 5'hd ? _GEN_1552 : _GEN_1447; // @[NulCtrlMP.scala 499:34]
  wire [4:0] _GEN_1697 = state == 5'hd ? _GEN_1682 : _GEN_1448; // @[NulCtrlMP.scala 499:34]
  wire [4:0] _GEN_1698 = state == 5'hd ? _GEN_1683 : _GEN_1449; // @[NulCtrlMP.scala 499:34]
  wire [4:0] _GEN_1699 = state == 5'hd ? _GEN_1684 : _GEN_1450; // @[NulCtrlMP.scala 499:34]
  wire [4:0] _GEN_1700 = state == 5'hd ? _GEN_1685 : _GEN_1451; // @[NulCtrlMP.scala 499:34]
  wire [128:0] _GEN_1701 = state == 5'hd ? _GEN_1691 : _GEN_1513; // @[NulCtrlMP.scala 499:34]
  wire [63:0] _GEN_1702 = state == 5'hd ? _GEN_1538 : _GEN_1453; // @[NulCtrlMP.scala 499:34]
  wire [63:0] _GEN_1703 = state == 5'hd ? _GEN_1558 : regback_1; // @[NulCtrlMP.scala 346:26 499:34]
  wire  _GEN_1704 = state == 5'hd ? _GEN_1678 : _GEN_1454; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1705 = state == 5'hd ? _GEN_1679 : _GEN_1455; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1706 = state == 5'hd ? _GEN_1680 : _GEN_1456; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1707 = state == 5'hd ? _GEN_1681 : _GEN_1457; // @[NulCtrlMP.scala 499:34]
  wire [63:0] _GEN_1708 = state == 5'hd ? _GEN_1686 : _GEN_1458; // @[NulCtrlMP.scala 499:34]
  wire [63:0] _GEN_1709 = state == 5'hd ? _GEN_1687 : _GEN_1459; // @[NulCtrlMP.scala 499:34]
  wire [63:0] _GEN_1710 = state == 5'hd ? _GEN_1688 : _GEN_1460; // @[NulCtrlMP.scala 499:34]
  wire [63:0] _GEN_1711 = state == 5'hd ? _GEN_1689 : _GEN_1461; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1712 = state == 5'hd ? _GEN_1620 : _GEN_1505; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1713 = state == 5'hd ? _GEN_1621 : _GEN_1506; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1714 = state == 5'hd ? _GEN_1622 : _GEN_1507; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1715 = state == 5'hd ? _GEN_1623 : _GEN_1508; // @[NulCtrlMP.scala 499:34]
  wire [31:0] _GEN_1716 = state == 5'hd ? _GEN_1624 : _GEN_1509; // @[NulCtrlMP.scala 499:34]
  wire [31:0] _GEN_1717 = state == 5'hd ? _GEN_1625 : _GEN_1510; // @[NulCtrlMP.scala 499:34]
  wire [31:0] _GEN_1718 = state == 5'hd ? _GEN_1626 : _GEN_1511; // @[NulCtrlMP.scala 499:34]
  wire [31:0] _GEN_1719 = state == 5'hd ? _GEN_1627 : _GEN_1512; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1720 = state == 5'hd ? _GEN_1634 : _GEN_1514; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1721 = state == 5'hd ? _GEN_1635 : _GEN_1515; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1722 = state == 5'hd ? _GEN_1636 : _GEN_1516; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1723 = state == 5'hd ? _GEN_1637 : _GEN_1517; // @[NulCtrlMP.scala 499:34]
  wire [4:0] _GEN_1724 = state == 5'hd ? _GEN_1692 : _GEN_1518; // @[NulCtrlMP.scala 499:34]
  wire  _GEN_1725 = _GEN_145 | _GEN_1712; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1726 = _GEN_146 | _GEN_1713; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1727 = _GEN_147 | _GEN_1714; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1728 = _GEN_148 | _GEN_1715; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_1729 = 2'h0 == opidx ? 32'h100f : _GEN_1716; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1730 = 2'h1 == opidx ? 32'h100f : _GEN_1717; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1731 = 2'h2 == opidx ? 32'h100f : _GEN_1718; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1732 = 2'h3 == opidx ? 32'h100f : _GEN_1719; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_1733 = _GEN_1180 ? _cnt_T : _GEN_1701; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1734 = cnt[0] ? _GEN_1725 : _GEN_1712; // @[NulCtrlMP.scala 513:22]
  wire  _GEN_1735 = cnt[0] ? _GEN_1726 : _GEN_1713; // @[NulCtrlMP.scala 513:22]
  wire  _GEN_1736 = cnt[0] ? _GEN_1727 : _GEN_1714; // @[NulCtrlMP.scala 513:22]
  wire  _GEN_1737 = cnt[0] ? _GEN_1728 : _GEN_1715; // @[NulCtrlMP.scala 513:22]
  wire [31:0] _GEN_1738 = cnt[0] ? _GEN_1729 : _GEN_1716; // @[NulCtrlMP.scala 513:22]
  wire [31:0] _GEN_1739 = cnt[0] ? _GEN_1730 : _GEN_1717; // @[NulCtrlMP.scala 513:22]
  wire [31:0] _GEN_1740 = cnt[0] ? _GEN_1731 : _GEN_1718; // @[NulCtrlMP.scala 513:22]
  wire [31:0] _GEN_1741 = cnt[0] ? _GEN_1732 : _GEN_1719; // @[NulCtrlMP.scala 513:22]
  wire [128:0] _GEN_1742 = cnt[0] ? _GEN_1733 : _GEN_1701; // @[NulCtrlMP.scala 513:22]
  wire  _GEN_1743 = _GEN_145 | _GEN_1720; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1744 = _GEN_146 | _GEN_1721; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1745 = _GEN_147 | _GEN_1722; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1746 = _GEN_148 | _GEN_1723; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_1747 = ~_GEN_1252 ? _cnt_T : _GEN_1742; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_1748 = cnt[1] ? _GEN_1743 : _GEN_1720; // @[NulCtrlMP.scala 514:22]
  wire  _GEN_1749 = cnt[1] ? _GEN_1744 : _GEN_1721; // @[NulCtrlMP.scala 514:22]
  wire  _GEN_1750 = cnt[1] ? _GEN_1745 : _GEN_1722; // @[NulCtrlMP.scala 514:22]
  wire  _GEN_1751 = cnt[1] ? _GEN_1746 : _GEN_1723; // @[NulCtrlMP.scala 514:22]
  wire [128:0] _GEN_1752 = cnt[1] ? _GEN_1747 : _GEN_1742; // @[NulCtrlMP.scala 514:22]
  wire [128:0] _GEN_1753 = cnt[2] ? 129'h1 : _GEN_1752; // @[NulCtrlMP.scala 515:22 516:17]
  wire [4:0] _GEN_1754 = cnt[2] ? 5'h5 : _GEN_1724; // @[NulCtrlMP.scala 515:22 517:19]
  wire  _GEN_1755 = state == 5'h16 ? _GEN_1734 : _GEN_1712; // @[NulCtrlMP.scala 512:33]
  wire  _GEN_1756 = state == 5'h16 ? _GEN_1735 : _GEN_1713; // @[NulCtrlMP.scala 512:33]
  wire  _GEN_1757 = state == 5'h16 ? _GEN_1736 : _GEN_1714; // @[NulCtrlMP.scala 512:33]
  wire  _GEN_1758 = state == 5'h16 ? _GEN_1737 : _GEN_1715; // @[NulCtrlMP.scala 512:33]
  wire [31:0] _GEN_1759 = state == 5'h16 ? _GEN_1738 : _GEN_1716; // @[NulCtrlMP.scala 512:33]
  wire [31:0] _GEN_1760 = state == 5'h16 ? _GEN_1739 : _GEN_1717; // @[NulCtrlMP.scala 512:33]
  wire [31:0] _GEN_1761 = state == 5'h16 ? _GEN_1740 : _GEN_1718; // @[NulCtrlMP.scala 512:33]
  wire [31:0] _GEN_1762 = state == 5'h16 ? _GEN_1741 : _GEN_1719; // @[NulCtrlMP.scala 512:33]
  wire [128:0] _GEN_1763 = state == 5'h16 ? _GEN_1753 : _GEN_1701; // @[NulCtrlMP.scala 512:33]
  wire  _GEN_1764 = state == 5'h16 ? _GEN_1748 : _GEN_1720; // @[NulCtrlMP.scala 512:33]
  wire  _GEN_1765 = state == 5'h16 ? _GEN_1749 : _GEN_1721; // @[NulCtrlMP.scala 512:33]
  wire  _GEN_1766 = state == 5'h16 ? _GEN_1750 : _GEN_1722; // @[NulCtrlMP.scala 512:33]
  wire  _GEN_1767 = state == 5'h16 ? _GEN_1751 : _GEN_1723; // @[NulCtrlMP.scala 512:33]
  wire [4:0] _GEN_1768 = state == 5'h16 ? _GEN_1754 : _GEN_1724; // @[NulCtrlMP.scala 512:33]
  wire  _T_181 = state == 5'he; // @[NulCtrlMP.scala 521:16]
  wire  _T_183 = ~oparg_2[5]; // @[NulCtrlMP.scala 521:35]
  wire  _GEN_1769 = _GEN_145 | _GEN_1693; // @[NulCtrlMP.scala 522:{27,27}]
  wire  _GEN_1770 = _GEN_146 | _GEN_1694; // @[NulCtrlMP.scala 522:{27,27}]
  wire  _GEN_1771 = _GEN_147 | _GEN_1695; // @[NulCtrlMP.scala 522:{27,27}]
  wire  _GEN_1772 = _GEN_148 | _GEN_1696; // @[NulCtrlMP.scala 522:{27,27}]
  wire [4:0] _GEN_1773 = 2'h0 == opidx ? oparg_2[4:0] : _GEN_1697; // @[NulCtrlMP.scala 523:{28,28}]
  wire [4:0] _GEN_1774 = 2'h1 == opidx ? oparg_2[4:0] : _GEN_1698; // @[NulCtrlMP.scala 523:{28,28}]
  wire [4:0] _GEN_1775 = 2'h2 == opidx ? oparg_2[4:0] : _GEN_1699; // @[NulCtrlMP.scala 523:{28,28}]
  wire [4:0] _GEN_1776 = 2'h3 == opidx ? oparg_2[4:0] : _GEN_1700; // @[NulCtrlMP.scala 523:{28,28}]
  wire [4:0] _GEN_1777 = _T_122 ? 5'h5 : _GEN_1768; // @[NulCtrlMP.scala 524:36 525:19]
  wire [7:0] _GEN_1778 = _T_122 ? _GEN_1349[7:0] : _GEN_1110; // @[NulCtrlMP.scala 524:36 527:27]
  wire [7:0] _GEN_1779 = _T_122 ? _GEN_1349[15:8] : _GEN_1033; // @[NulCtrlMP.scala 524:36 527:27]
  wire [7:0] _GEN_1780 = _T_122 ? _GEN_1349[23:16] : _GEN_1034; // @[NulCtrlMP.scala 524:36 527:27]
  wire [7:0] _GEN_1781 = _T_122 ? _GEN_1349[31:24] : _GEN_1035; // @[NulCtrlMP.scala 524:36 527:27]
  wire [7:0] _GEN_1782 = _T_122 ? _GEN_1349[39:32] : _GEN_1036; // @[NulCtrlMP.scala 524:36 527:27]
  wire [7:0] _GEN_1783 = _T_122 ? _GEN_1349[47:40] : _GEN_1037; // @[NulCtrlMP.scala 524:36 527:27]
  wire [7:0] _GEN_1784 = _T_122 ? _GEN_1349[55:48] : _GEN_1038; // @[NulCtrlMP.scala 524:36 527:27]
  wire [7:0] _GEN_1785 = _T_122 ? _GEN_1349[63:56] : _GEN_1039; // @[NulCtrlMP.scala 524:36 527:27]
  wire  _GEN_1786 = state == 5'he & ~oparg_2[5] ? _GEN_1769 : _GEN_1693; // @[NulCtrlMP.scala 521:49]
  wire  _GEN_1787 = state == 5'he & ~oparg_2[5] ? _GEN_1770 : _GEN_1694; // @[NulCtrlMP.scala 521:49]
  wire  _GEN_1788 = state == 5'he & ~oparg_2[5] ? _GEN_1771 : _GEN_1695; // @[NulCtrlMP.scala 521:49]
  wire  _GEN_1789 = state == 5'he & ~oparg_2[5] ? _GEN_1772 : _GEN_1696; // @[NulCtrlMP.scala 521:49]
  wire [4:0] _GEN_1790 = state == 5'he & ~oparg_2[5] ? _GEN_1773 : _GEN_1697; // @[NulCtrlMP.scala 521:49]
  wire [4:0] _GEN_1791 = state == 5'he & ~oparg_2[5] ? _GEN_1774 : _GEN_1698; // @[NulCtrlMP.scala 521:49]
  wire [4:0] _GEN_1792 = state == 5'he & ~oparg_2[5] ? _GEN_1775 : _GEN_1699; // @[NulCtrlMP.scala 521:49]
  wire [4:0] _GEN_1793 = state == 5'he & ~oparg_2[5] ? _GEN_1776 : _GEN_1700; // @[NulCtrlMP.scala 521:49]
  wire [4:0] _GEN_1794 = state == 5'he & ~oparg_2[5] ? _GEN_1777 : _GEN_1768; // @[NulCtrlMP.scala 521:49]
  wire [7:0] _GEN_1795 = state == 5'he & ~oparg_2[5] ? _GEN_1778 : _GEN_1110; // @[NulCtrlMP.scala 521:49]
  wire [7:0] _GEN_1796 = state == 5'he & ~oparg_2[5] ? _GEN_1779 : _GEN_1033; // @[NulCtrlMP.scala 521:49]
  wire [7:0] _GEN_1797 = state == 5'he & ~oparg_2[5] ? _GEN_1780 : _GEN_1034; // @[NulCtrlMP.scala 521:49]
  wire [7:0] _GEN_1798 = state == 5'he & ~oparg_2[5] ? _GEN_1781 : _GEN_1035; // @[NulCtrlMP.scala 521:49]
  wire [7:0] _GEN_1799 = state == 5'he & ~oparg_2[5] ? _GEN_1782 : _GEN_1036; // @[NulCtrlMP.scala 521:49]
  wire [7:0] _GEN_1800 = state == 5'he & ~oparg_2[5] ? _GEN_1783 : _GEN_1037; // @[NulCtrlMP.scala 521:49]
  wire [7:0] _GEN_1801 = state == 5'he & ~oparg_2[5] ? _GEN_1784 : _GEN_1038; // @[NulCtrlMP.scala 521:49]
  wire [7:0] _GEN_1802 = state == 5'he & ~oparg_2[5] ? _GEN_1785 : _GEN_1039; // @[NulCtrlMP.scala 521:49]
  wire  _GEN_1803 = _GEN_145 | _GEN_1786; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1804 = _GEN_146 | _GEN_1787; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1805 = _GEN_147 | _GEN_1788; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1806 = _GEN_148 | _GEN_1789; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_1807 = 2'h0 == opidx ? 5'h5 : _GEN_1790; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1808 = 2'h1 == opidx ? 5'h5 : _GEN_1791; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1809 = 2'h2 == opidx ? 5'h5 : _GEN_1792; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1810 = 2'h3 == opidx ? 5'h5 : _GEN_1793; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_1811 = _T_122 ? _cnt_T : _GEN_1763; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_1812 = _T_122 ? _GEN_1349 : _GEN_1702; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_1813 = cnt[0] ? _GEN_1803 : _GEN_1786; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1814 = cnt[0] ? _GEN_1804 : _GEN_1787; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1815 = cnt[0] ? _GEN_1805 : _GEN_1788; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1816 = cnt[0] ? _GEN_1806 : _GEN_1789; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1817 = cnt[0] ? _GEN_1807 : _GEN_1790; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1818 = cnt[0] ? _GEN_1808 : _GEN_1791; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1819 = cnt[0] ? _GEN_1809 : _GEN_1792; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1820 = cnt[0] ? _GEN_1810 : _GEN_1793; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_1821 = cnt[0] ? _GEN_1811 : _GEN_1763; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_1822 = cnt[0] ? _GEN_1812 : _GEN_1702; // @[NulCtrlMP.scala 408:32]
  wire [19:0] _T_193 = {oparg_2[4:0], 15'h0}; // @[NulCtrlMP.scala 534:70]
  wire [31:0] _GEN_9290 = {{12'd0}, _T_193}; // @[NulCtrlMP.scala 534:52]
  wire [31:0] _T_194 = 32'he20002d3 | _GEN_9290; // @[NulCtrlMP.scala 534:52]
  wire  _GEN_1823 = _GEN_145 | _GEN_1755; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1824 = _GEN_146 | _GEN_1756; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1825 = _GEN_147 | _GEN_1757; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_1826 = _GEN_148 | _GEN_1758; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_1827 = 2'h0 == opidx ? _T_194 : _GEN_1759; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1828 = 2'h1 == opidx ? _T_194 : _GEN_1760; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1829 = 2'h2 == opidx ? _T_194 : _GEN_1761; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_1830 = 2'h3 == opidx ? _T_194 : _GEN_1762; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_1831 = _GEN_1180 ? _cnt_T : _GEN_1821; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_1832 = cnt[1] ? _GEN_1823 : _GEN_1755; // @[NulCtrlMP.scala 534:22]
  wire  _GEN_1833 = cnt[1] ? _GEN_1824 : _GEN_1756; // @[NulCtrlMP.scala 534:22]
  wire  _GEN_1834 = cnt[1] ? _GEN_1825 : _GEN_1757; // @[NulCtrlMP.scala 534:22]
  wire  _GEN_1835 = cnt[1] ? _GEN_1826 : _GEN_1758; // @[NulCtrlMP.scala 534:22]
  wire [31:0] _GEN_1836 = cnt[1] ? _GEN_1827 : _GEN_1759; // @[NulCtrlMP.scala 534:22]
  wire [31:0] _GEN_1837 = cnt[1] ? _GEN_1828 : _GEN_1760; // @[NulCtrlMP.scala 534:22]
  wire [31:0] _GEN_1838 = cnt[1] ? _GEN_1829 : _GEN_1761; // @[NulCtrlMP.scala 534:22]
  wire [31:0] _GEN_1839 = cnt[1] ? _GEN_1830 : _GEN_1762; // @[NulCtrlMP.scala 534:22]
  wire [128:0] _GEN_1840 = cnt[1] ? _GEN_1831 : _GEN_1821; // @[NulCtrlMP.scala 534:22]
  wire  _GEN_1841 = _GEN_145 | _GEN_1764; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1842 = _GEN_146 | _GEN_1765; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1843 = _GEN_147 | _GEN_1766; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_1844 = _GEN_148 | _GEN_1767; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_1845 = ~_GEN_1252 ? _cnt_T : _GEN_1840; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_1846 = cnt[2] ? _GEN_1841 : _GEN_1764; // @[NulCtrlMP.scala 535:22]
  wire  _GEN_1847 = cnt[2] ? _GEN_1842 : _GEN_1765; // @[NulCtrlMP.scala 535:22]
  wire  _GEN_1848 = cnt[2] ? _GEN_1843 : _GEN_1766; // @[NulCtrlMP.scala 535:22]
  wire  _GEN_1849 = cnt[2] ? _GEN_1844 : _GEN_1767; // @[NulCtrlMP.scala 535:22]
  wire [128:0] _GEN_1850 = cnt[2] ? _GEN_1845 : _GEN_1840; // @[NulCtrlMP.scala 535:22]
  wire  _GEN_1851 = _GEN_145 | _GEN_1813; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_1852 = _GEN_146 | _GEN_1814; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_1853 = _GEN_147 | _GEN_1815; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_1854 = _GEN_148 | _GEN_1816; // @[NulCtrlMP.scala 359:{27,27}]
  wire [4:0] _GEN_1855 = 2'h0 == opidx ? 5'h5 : _GEN_1817; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_1856 = 2'h1 == opidx ? 5'h5 : _GEN_1818; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_1857 = 2'h2 == opidx ? 5'h5 : _GEN_1819; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_1858 = 2'h3 == opidx ? 5'h5 : _GEN_1820; // @[NulCtrlMP.scala 360:{28,28}]
  wire [128:0] _GEN_1859 = _T_122 ? _cnt_T : _GEN_1850; // @[NulCtrlMP.scala 361:36 362:17]
  wire [7:0] _GEN_1860 = _T_122 ? _GEN_1349[7:0] : _GEN_1797; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_1861 = _T_122 ? _GEN_1349[15:8] : _GEN_1798; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_1862 = _T_122 ? _GEN_1349[23:16] : _GEN_1799; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_1863 = _T_122 ? _GEN_1349[31:24] : _GEN_1800; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_1864 = _T_122 ? _GEN_1349[39:32] : _GEN_1801; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_1865 = _T_122 ? _GEN_1349[47:40] : _GEN_1802; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_1866 = _T_122 ? _GEN_1349[55:48] : retarg_8; // @[NulCtrlMP.scala 152:25 361:36 364:33]
  wire [7:0] _GEN_1867 = _T_122 ? _GEN_1349[63:56] : retarg_9; // @[NulCtrlMP.scala 152:25 361:36 364:33]
  wire  _GEN_1868 = cnt[3] ? _GEN_1851 : _GEN_1813; // @[NulCtrlMP.scala 536:22]
  wire  _GEN_1869 = cnt[3] ? _GEN_1852 : _GEN_1814; // @[NulCtrlMP.scala 536:22]
  wire  _GEN_1870 = cnt[3] ? _GEN_1853 : _GEN_1815; // @[NulCtrlMP.scala 536:22]
  wire  _GEN_1871 = cnt[3] ? _GEN_1854 : _GEN_1816; // @[NulCtrlMP.scala 536:22]
  wire [4:0] _GEN_1872 = cnt[3] ? _GEN_1855 : _GEN_1817; // @[NulCtrlMP.scala 536:22]
  wire [4:0] _GEN_1873 = cnt[3] ? _GEN_1856 : _GEN_1818; // @[NulCtrlMP.scala 536:22]
  wire [4:0] _GEN_1874 = cnt[3] ? _GEN_1857 : _GEN_1819; // @[NulCtrlMP.scala 536:22]
  wire [4:0] _GEN_1875 = cnt[3] ? _GEN_1858 : _GEN_1820; // @[NulCtrlMP.scala 536:22]
  wire [128:0] _GEN_1876 = cnt[3] ? _GEN_1859 : _GEN_1850; // @[NulCtrlMP.scala 536:22]
  wire [7:0] _GEN_1877 = cnt[3] ? _GEN_1860 : _GEN_1797; // @[NulCtrlMP.scala 536:22]
  wire [7:0] _GEN_1878 = cnt[3] ? _GEN_1861 : _GEN_1798; // @[NulCtrlMP.scala 536:22]
  wire [7:0] _GEN_1879 = cnt[3] ? _GEN_1862 : _GEN_1799; // @[NulCtrlMP.scala 536:22]
  wire [7:0] _GEN_1880 = cnt[3] ? _GEN_1863 : _GEN_1800; // @[NulCtrlMP.scala 536:22]
  wire [7:0] _GEN_1881 = cnt[3] ? _GEN_1864 : _GEN_1801; // @[NulCtrlMP.scala 536:22]
  wire [7:0] _GEN_1882 = cnt[3] ? _GEN_1865 : _GEN_1802; // @[NulCtrlMP.scala 536:22]
  wire [7:0] _GEN_1883 = cnt[3] ? _GEN_1866 : retarg_8; // @[NulCtrlMP.scala 536:22 152:25]
  wire [7:0] _GEN_1884 = cnt[3] ? _GEN_1867 : retarg_9; // @[NulCtrlMP.scala 536:22 152:25]
  wire  _GEN_1885 = _GEN_145 | _GEN_1704; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1886 = _GEN_146 | _GEN_1705; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1887 = _GEN_147 | _GEN_1706; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_1888 = _GEN_148 | _GEN_1707; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_1889 = 2'h0 == opidx ? 5'h5 : _GEN_1872; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1890 = 2'h1 == opidx ? 5'h5 : _GEN_1873; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1891 = 2'h2 == opidx ? 5'h5 : _GEN_1874; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_1892 = 2'h3 == opidx ? 5'h5 : _GEN_1875; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_1893 = 2'h0 == opidx ? regback_0 : _GEN_1708; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1894 = 2'h1 == opidx ? regback_0 : _GEN_1709; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1895 = 2'h2 == opidx ? regback_0 : _GEN_1710; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_1896 = 2'h3 == opidx ? regback_0 : _GEN_1711; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_1897 = ~_GEN_1128 ? _cnt_T : _GEN_1876; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_1898 = cnt[4] ? _GEN_1885 : _GEN_1704; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1899 = cnt[4] ? _GEN_1886 : _GEN_1705; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1900 = cnt[4] ? _GEN_1887 : _GEN_1706; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_1901 = cnt[4] ? _GEN_1888 : _GEN_1707; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1902 = cnt[4] ? _GEN_1889 : _GEN_1872; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1903 = cnt[4] ? _GEN_1890 : _GEN_1873; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1904 = cnt[4] ? _GEN_1891 : _GEN_1874; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_1905 = cnt[4] ? _GEN_1892 : _GEN_1875; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1906 = cnt[4] ? _GEN_1893 : _GEN_1708; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1907 = cnt[4] ? _GEN_1894 : _GEN_1709; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1908 = cnt[4] ? _GEN_1895 : _GEN_1710; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_1909 = cnt[4] ? _GEN_1896 : _GEN_1711; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_1910 = cnt[4] ? _GEN_1897 : _GEN_1876; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_1911 = cnt[5] ? 129'h1 : _GEN_1910; // @[NulCtrlMP.scala 538:22 539:17]
  wire [4:0] _GEN_1912 = cnt[5] ? 5'h5 : _GEN_1794; // @[NulCtrlMP.scala 538:22 540:19]
  wire  _GEN_1913 = _T_181 & oparg_2[5] ? _GEN_1868 : _GEN_1786; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1914 = _T_181 & oparg_2[5] ? _GEN_1869 : _GEN_1787; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1915 = _T_181 & oparg_2[5] ? _GEN_1870 : _GEN_1788; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1916 = _T_181 & oparg_2[5] ? _GEN_1871 : _GEN_1789; // @[NulCtrlMP.scala 532:48]
  wire [4:0] _GEN_1917 = _T_181 & oparg_2[5] ? _GEN_1902 : _GEN_1790; // @[NulCtrlMP.scala 532:48]
  wire [4:0] _GEN_1918 = _T_181 & oparg_2[5] ? _GEN_1903 : _GEN_1791; // @[NulCtrlMP.scala 532:48]
  wire [4:0] _GEN_1919 = _T_181 & oparg_2[5] ? _GEN_1904 : _GEN_1792; // @[NulCtrlMP.scala 532:48]
  wire [4:0] _GEN_1920 = _T_181 & oparg_2[5] ? _GEN_1905 : _GEN_1793; // @[NulCtrlMP.scala 532:48]
  wire [128:0] _GEN_1921 = _T_181 & oparg_2[5] ? _GEN_1911 : _GEN_1763; // @[NulCtrlMP.scala 532:48]
  wire [63:0] _GEN_1922 = _T_181 & oparg_2[5] ? _GEN_1822 : _GEN_1702; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1923 = _T_181 & oparg_2[5] ? _GEN_1832 : _GEN_1755; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1924 = _T_181 & oparg_2[5] ? _GEN_1833 : _GEN_1756; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1925 = _T_181 & oparg_2[5] ? _GEN_1834 : _GEN_1757; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1926 = _T_181 & oparg_2[5] ? _GEN_1835 : _GEN_1758; // @[NulCtrlMP.scala 532:48]
  wire [31:0] _GEN_1927 = _T_181 & oparg_2[5] ? _GEN_1836 : _GEN_1759; // @[NulCtrlMP.scala 532:48]
  wire [31:0] _GEN_1928 = _T_181 & oparg_2[5] ? _GEN_1837 : _GEN_1760; // @[NulCtrlMP.scala 532:48]
  wire [31:0] _GEN_1929 = _T_181 & oparg_2[5] ? _GEN_1838 : _GEN_1761; // @[NulCtrlMP.scala 532:48]
  wire [31:0] _GEN_1930 = _T_181 & oparg_2[5] ? _GEN_1839 : _GEN_1762; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1931 = _T_181 & oparg_2[5] ? _GEN_1846 : _GEN_1764; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1932 = _T_181 & oparg_2[5] ? _GEN_1847 : _GEN_1765; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1933 = _T_181 & oparg_2[5] ? _GEN_1848 : _GEN_1766; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1934 = _T_181 & oparg_2[5] ? _GEN_1849 : _GEN_1767; // @[NulCtrlMP.scala 532:48]
  wire [7:0] _GEN_1935 = _T_181 & oparg_2[5] ? _GEN_1877 : _GEN_1797; // @[NulCtrlMP.scala 532:48]
  wire [7:0] _GEN_1936 = _T_181 & oparg_2[5] ? _GEN_1878 : _GEN_1798; // @[NulCtrlMP.scala 532:48]
  wire [7:0] _GEN_1937 = _T_181 & oparg_2[5] ? _GEN_1879 : _GEN_1799; // @[NulCtrlMP.scala 532:48]
  wire [7:0] _GEN_1938 = _T_181 & oparg_2[5] ? _GEN_1880 : _GEN_1800; // @[NulCtrlMP.scala 532:48]
  wire [7:0] _GEN_1939 = _T_181 & oparg_2[5] ? _GEN_1881 : _GEN_1801; // @[NulCtrlMP.scala 532:48]
  wire [7:0] _GEN_1940 = _T_181 & oparg_2[5] ? _GEN_1882 : _GEN_1802; // @[NulCtrlMP.scala 532:48]
  wire [7:0] _GEN_1941 = _T_181 & oparg_2[5] ? _GEN_1883 : retarg_8; // @[NulCtrlMP.scala 152:25 532:48]
  wire [7:0] _GEN_1942 = _T_181 & oparg_2[5] ? _GEN_1884 : retarg_9; // @[NulCtrlMP.scala 152:25 532:48]
  wire  _GEN_1943 = _T_181 & oparg_2[5] ? _GEN_1898 : _GEN_1704; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1944 = _T_181 & oparg_2[5] ? _GEN_1899 : _GEN_1705; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1945 = _T_181 & oparg_2[5] ? _GEN_1900 : _GEN_1706; // @[NulCtrlMP.scala 532:48]
  wire  _GEN_1946 = _T_181 & oparg_2[5] ? _GEN_1901 : _GEN_1707; // @[NulCtrlMP.scala 532:48]
  wire [63:0] _GEN_1947 = _T_181 & oparg_2[5] ? _GEN_1906 : _GEN_1708; // @[NulCtrlMP.scala 532:48]
  wire [63:0] _GEN_1948 = _T_181 & oparg_2[5] ? _GEN_1907 : _GEN_1709; // @[NulCtrlMP.scala 532:48]
  wire [63:0] _GEN_1949 = _T_181 & oparg_2[5] ? _GEN_1908 : _GEN_1710; // @[NulCtrlMP.scala 532:48]
  wire [63:0] _GEN_1950 = _T_181 & oparg_2[5] ? _GEN_1909 : _GEN_1711; // @[NulCtrlMP.scala 532:48]
  wire [4:0] _GEN_1951 = _T_181 & oparg_2[5] ? _GEN_1912 : _GEN_1794; // @[NulCtrlMP.scala 532:48]
  wire  _T_202 = state == 5'hf; // @[NulCtrlMP.scala 544:16]
  wire  _GEN_1952 = _GEN_145 | _GEN_1943; // @[NulCtrlMP.scala 545:{27,27}]
  wire  _GEN_1953 = _GEN_146 | _GEN_1944; // @[NulCtrlMP.scala 545:{27,27}]
  wire  _GEN_1954 = _GEN_147 | _GEN_1945; // @[NulCtrlMP.scala 545:{27,27}]
  wire  _GEN_1955 = _GEN_148 | _GEN_1946; // @[NulCtrlMP.scala 545:{27,27}]
  wire [4:0] _GEN_1956 = 2'h0 == opidx ? oparg_2[4:0] : _GEN_1917; // @[NulCtrlMP.scala 546:{28,28}]
  wire [4:0] _GEN_1957 = 2'h1 == opidx ? oparg_2[4:0] : _GEN_1918; // @[NulCtrlMP.scala 546:{28,28}]
  wire [4:0] _GEN_1958 = 2'h2 == opidx ? oparg_2[4:0] : _GEN_1919; // @[NulCtrlMP.scala 546:{28,28}]
  wire [4:0] _GEN_1959 = 2'h3 == opidx ? oparg_2[4:0] : _GEN_1920; // @[NulCtrlMP.scala 546:{28,28}]
  wire [63:0] _io_cpu_regacc_wdata_T = {oparg_11,oparg_10,oparg_9,oparg_8,oparg_7,oparg_6,oparg_5,oparg_4}; // @[NulCtrlMP.scala 551:53]
  wire [63:0] _GEN_1960 = 2'h0 == opidx ? _io_cpu_regacc_wdata_T : _GEN_1947; // @[NulCtrlMP.scala 551:{30,30}]
  wire [63:0] _GEN_1961 = 2'h1 == opidx ? _io_cpu_regacc_wdata_T : _GEN_1948; // @[NulCtrlMP.scala 551:{30,30}]
  wire [63:0] _GEN_1962 = 2'h2 == opidx ? _io_cpu_regacc_wdata_T : _GEN_1949; // @[NulCtrlMP.scala 551:{30,30}]
  wire [63:0] _GEN_1963 = 2'h3 == opidx ? _io_cpu_regacc_wdata_T : _GEN_1950; // @[NulCtrlMP.scala 551:{30,30}]
  wire [4:0] _GEN_1964 = _T_122 ? 5'h5 : _GEN_1951; // @[NulCtrlMP.scala 552:36 553:19]
  wire  _GEN_1965 = state == 5'hf & _T_183 ? _GEN_1952 : _GEN_1943; // @[NulCtrlMP.scala 544:49]
  wire  _GEN_1966 = state == 5'hf & _T_183 ? _GEN_1953 : _GEN_1944; // @[NulCtrlMP.scala 544:49]
  wire  _GEN_1967 = state == 5'hf & _T_183 ? _GEN_1954 : _GEN_1945; // @[NulCtrlMP.scala 544:49]
  wire  _GEN_1968 = state == 5'hf & _T_183 ? _GEN_1955 : _GEN_1946; // @[NulCtrlMP.scala 544:49]
  wire [4:0] _GEN_1969 = state == 5'hf & _T_183 ? _GEN_1956 : _GEN_1917; // @[NulCtrlMP.scala 544:49]
  wire [4:0] _GEN_1970 = state == 5'hf & _T_183 ? _GEN_1957 : _GEN_1918; // @[NulCtrlMP.scala 544:49]
  wire [4:0] _GEN_1971 = state == 5'hf & _T_183 ? _GEN_1958 : _GEN_1919; // @[NulCtrlMP.scala 544:49]
  wire [4:0] _GEN_1972 = state == 5'hf & _T_183 ? _GEN_1959 : _GEN_1920; // @[NulCtrlMP.scala 544:49]
  wire [63:0] _GEN_1973 = state == 5'hf & _T_183 ? _GEN_1960 : _GEN_1947; // @[NulCtrlMP.scala 544:49]
  wire [63:0] _GEN_1974 = state == 5'hf & _T_183 ? _GEN_1961 : _GEN_1948; // @[NulCtrlMP.scala 544:49]
  wire [63:0] _GEN_1975 = state == 5'hf & _T_183 ? _GEN_1962 : _GEN_1949; // @[NulCtrlMP.scala 544:49]
  wire [63:0] _GEN_1976 = state == 5'hf & _T_183 ? _GEN_1963 : _GEN_1950; // @[NulCtrlMP.scala 544:49]
  wire [4:0] _GEN_1977 = state == 5'hf & _T_183 ? _GEN_1964 : _GEN_1951; // @[NulCtrlMP.scala 544:49]
  wire  _GEN_1978 = _GEN_145 | _GEN_1913; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1979 = _GEN_146 | _GEN_1914; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1980 = _GEN_147 | _GEN_1915; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_1981 = _GEN_148 | _GEN_1916; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_1982 = 2'h0 == opidx ? 5'h5 : _GEN_1969; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1983 = 2'h1 == opidx ? 5'h5 : _GEN_1970; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1984 = 2'h2 == opidx ? 5'h5 : _GEN_1971; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_1985 = 2'h3 == opidx ? 5'h5 : _GEN_1972; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_1986 = _T_122 ? _cnt_T : _GEN_1921; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_1987 = _T_122 ? _GEN_1349 : _GEN_1922; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_1988 = cnt[0] ? _GEN_1978 : _GEN_1913; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1989 = cnt[0] ? _GEN_1979 : _GEN_1914; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1990 = cnt[0] ? _GEN_1980 : _GEN_1915; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1991 = cnt[0] ? _GEN_1981 : _GEN_1916; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1992 = cnt[0] ? _GEN_1982 : _GEN_1969; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1993 = cnt[0] ? _GEN_1983 : _GEN_1970; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1994 = cnt[0] ? _GEN_1984 : _GEN_1971; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_1995 = cnt[0] ? _GEN_1985 : _GEN_1972; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_1996 = cnt[0] ? _GEN_1986 : _GEN_1921; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_1997 = cnt[0] ? _GEN_1987 : _GEN_1922; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_1998 = _GEN_145 | _GEN_1965; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_1999 = _GEN_146 | _GEN_1966; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_2000 = _GEN_147 | _GEN_1967; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_2001 = _GEN_148 | _GEN_1968; // @[NulCtrlMP.scala 377:{27,27}]
  wire [4:0] _GEN_2002 = 2'h0 == opidx ? 5'h5 : _GEN_1992; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_2003 = 2'h1 == opidx ? 5'h5 : _GEN_1993; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_2004 = 2'h2 == opidx ? 5'h5 : _GEN_1994; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_2005 = 2'h3 == opidx ? 5'h5 : _GEN_1995; // @[NulCtrlMP.scala 378:{28,28}]
  wire [63:0] _GEN_2006 = 2'h0 == opidx ? _io_cpu_regacc_wdata_T : _GEN_1973; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_2007 = 2'h1 == opidx ? _io_cpu_regacc_wdata_T : _GEN_1974; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_2008 = 2'h2 == opidx ? _io_cpu_regacc_wdata_T : _GEN_1975; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_2009 = 2'h3 == opidx ? _io_cpu_regacc_wdata_T : _GEN_1976; // @[NulCtrlMP.scala 388:{30,30}]
  wire [128:0] _GEN_2010 = _T_122 ? _cnt_T : _GEN_1996; // @[NulCtrlMP.scala 389:36 390:17]
  wire  _GEN_2011 = cnt[1] ? _GEN_1998 : _GEN_1965; // @[NulCtrlMP.scala 559:22]
  wire  _GEN_2012 = cnt[1] ? _GEN_1999 : _GEN_1966; // @[NulCtrlMP.scala 559:22]
  wire  _GEN_2013 = cnt[1] ? _GEN_2000 : _GEN_1967; // @[NulCtrlMP.scala 559:22]
  wire  _GEN_2014 = cnt[1] ? _GEN_2001 : _GEN_1968; // @[NulCtrlMP.scala 559:22]
  wire [4:0] _GEN_2015 = cnt[1] ? _GEN_2002 : _GEN_1992; // @[NulCtrlMP.scala 559:22]
  wire [4:0] _GEN_2016 = cnt[1] ? _GEN_2003 : _GEN_1993; // @[NulCtrlMP.scala 559:22]
  wire [4:0] _GEN_2017 = cnt[1] ? _GEN_2004 : _GEN_1994; // @[NulCtrlMP.scala 559:22]
  wire [4:0] _GEN_2018 = cnt[1] ? _GEN_2005 : _GEN_1995; // @[NulCtrlMP.scala 559:22]
  wire [63:0] _GEN_2019 = cnt[1] ? _GEN_2006 : _GEN_1973; // @[NulCtrlMP.scala 559:22]
  wire [63:0] _GEN_2020 = cnt[1] ? _GEN_2007 : _GEN_1974; // @[NulCtrlMP.scala 559:22]
  wire [63:0] _GEN_2021 = cnt[1] ? _GEN_2008 : _GEN_1975; // @[NulCtrlMP.scala 559:22]
  wire [63:0] _GEN_2022 = cnt[1] ? _GEN_2009 : _GEN_1976; // @[NulCtrlMP.scala 559:22]
  wire [128:0] _GEN_2023 = cnt[1] ? _GEN_2010 : _GEN_1996; // @[NulCtrlMP.scala 559:22]
  wire [11:0] _T_216 = {oparg_2[4:0], 7'h0}; // @[NulCtrlMP.scala 560:70]
  wire [31:0] _GEN_9319 = {{20'd0}, _T_216}; // @[NulCtrlMP.scala 560:52]
  wire [31:0] _T_217 = 32'hf2028053 | _GEN_9319; // @[NulCtrlMP.scala 560:52]
  wire  _GEN_2024 = _GEN_145 | _GEN_1923; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2025 = _GEN_146 | _GEN_1924; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2026 = _GEN_147 | _GEN_1925; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2027 = _GEN_148 | _GEN_1926; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2028 = 2'h0 == opidx ? _T_217 : _GEN_1927; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2029 = 2'h1 == opidx ? _T_217 : _GEN_1928; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2030 = 2'h2 == opidx ? _T_217 : _GEN_1929; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2031 = 2'h3 == opidx ? _T_217 : _GEN_1930; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2032 = _GEN_1180 ? _cnt_T : _GEN_2023; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2033 = cnt[2] ? _GEN_2024 : _GEN_1923; // @[NulCtrlMP.scala 560:22]
  wire  _GEN_2034 = cnt[2] ? _GEN_2025 : _GEN_1924; // @[NulCtrlMP.scala 560:22]
  wire  _GEN_2035 = cnt[2] ? _GEN_2026 : _GEN_1925; // @[NulCtrlMP.scala 560:22]
  wire  _GEN_2036 = cnt[2] ? _GEN_2027 : _GEN_1926; // @[NulCtrlMP.scala 560:22]
  wire [31:0] _GEN_2037 = cnt[2] ? _GEN_2028 : _GEN_1927; // @[NulCtrlMP.scala 560:22]
  wire [31:0] _GEN_2038 = cnt[2] ? _GEN_2029 : _GEN_1928; // @[NulCtrlMP.scala 560:22]
  wire [31:0] _GEN_2039 = cnt[2] ? _GEN_2030 : _GEN_1929; // @[NulCtrlMP.scala 560:22]
  wire [31:0] _GEN_2040 = cnt[2] ? _GEN_2031 : _GEN_1930; // @[NulCtrlMP.scala 560:22]
  wire [128:0] _GEN_2041 = cnt[2] ? _GEN_2032 : _GEN_2023; // @[NulCtrlMP.scala 560:22]
  wire  _GEN_2042 = _GEN_145 | _GEN_1931; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_2043 = _GEN_146 | _GEN_1932; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_2044 = _GEN_147 | _GEN_1933; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_2045 = _GEN_148 | _GEN_1934; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_2046 = ~_GEN_1252 ? _cnt_T : _GEN_2041; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_2047 = cnt[3] ? _GEN_2042 : _GEN_1931; // @[NulCtrlMP.scala 561:22]
  wire  _GEN_2048 = cnt[3] ? _GEN_2043 : _GEN_1932; // @[NulCtrlMP.scala 561:22]
  wire  _GEN_2049 = cnt[3] ? _GEN_2044 : _GEN_1933; // @[NulCtrlMP.scala 561:22]
  wire  _GEN_2050 = cnt[3] ? _GEN_2045 : _GEN_1934; // @[NulCtrlMP.scala 561:22]
  wire [128:0] _GEN_2051 = cnt[3] ? _GEN_2046 : _GEN_2041; // @[NulCtrlMP.scala 561:22]
  wire  _GEN_2052 = _GEN_145 | _GEN_2011; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2053 = _GEN_146 | _GEN_2012; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2054 = _GEN_147 | _GEN_2013; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2055 = _GEN_148 | _GEN_2014; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_2056 = 2'h0 == opidx ? 5'h5 : _GEN_2015; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2057 = 2'h1 == opidx ? 5'h5 : _GEN_2016; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2058 = 2'h2 == opidx ? 5'h5 : _GEN_2017; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2059 = 2'h3 == opidx ? 5'h5 : _GEN_2018; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_2060 = 2'h0 == opidx ? regback_0 : _GEN_2019; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2061 = 2'h1 == opidx ? regback_0 : _GEN_2020; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2062 = 2'h2 == opidx ? regback_0 : _GEN_2021; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2063 = 2'h3 == opidx ? regback_0 : _GEN_2022; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_2064 = ~_GEN_1128 ? _cnt_T : _GEN_2051; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_2065 = cnt[4] ? _GEN_2052 : _GEN_2011; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2066 = cnt[4] ? _GEN_2053 : _GEN_2012; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2067 = cnt[4] ? _GEN_2054 : _GEN_2013; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2068 = cnt[4] ? _GEN_2055 : _GEN_2014; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2069 = cnt[4] ? _GEN_2056 : _GEN_2015; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2070 = cnt[4] ? _GEN_2057 : _GEN_2016; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2071 = cnt[4] ? _GEN_2058 : _GEN_2017; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2072 = cnt[4] ? _GEN_2059 : _GEN_2018; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2073 = cnt[4] ? _GEN_2060 : _GEN_2019; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2074 = cnt[4] ? _GEN_2061 : _GEN_2020; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2075 = cnt[4] ? _GEN_2062 : _GEN_2021; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2076 = cnt[4] ? _GEN_2063 : _GEN_2022; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_2077 = cnt[4] ? _GEN_2064 : _GEN_2051; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_2078 = cnt[5] ? 129'h1 : _GEN_2077; // @[NulCtrlMP.scala 563:22 564:17]
  wire [4:0] _GEN_2079 = cnt[5] ? 5'h5 : _GEN_1977; // @[NulCtrlMP.scala 563:22 565:19]
  wire  _GEN_2080 = _T_202 & oparg_2[5] ? _GEN_1988 : _GEN_1913; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2081 = _T_202 & oparg_2[5] ? _GEN_1989 : _GEN_1914; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2082 = _T_202 & oparg_2[5] ? _GEN_1990 : _GEN_1915; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2083 = _T_202 & oparg_2[5] ? _GEN_1991 : _GEN_1916; // @[NulCtrlMP.scala 557:48]
  wire [4:0] _GEN_2084 = _T_202 & oparg_2[5] ? _GEN_2069 : _GEN_1969; // @[NulCtrlMP.scala 557:48]
  wire [4:0] _GEN_2085 = _T_202 & oparg_2[5] ? _GEN_2070 : _GEN_1970; // @[NulCtrlMP.scala 557:48]
  wire [4:0] _GEN_2086 = _T_202 & oparg_2[5] ? _GEN_2071 : _GEN_1971; // @[NulCtrlMP.scala 557:48]
  wire [4:0] _GEN_2087 = _T_202 & oparg_2[5] ? _GEN_2072 : _GEN_1972; // @[NulCtrlMP.scala 557:48]
  wire [128:0] _GEN_2088 = _T_202 & oparg_2[5] ? _GEN_2078 : _GEN_1921; // @[NulCtrlMP.scala 557:48]
  wire [63:0] _GEN_2089 = _T_202 & oparg_2[5] ? _GEN_1997 : _GEN_1922; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2090 = _T_202 & oparg_2[5] ? _GEN_2065 : _GEN_1965; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2091 = _T_202 & oparg_2[5] ? _GEN_2066 : _GEN_1966; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2092 = _T_202 & oparg_2[5] ? _GEN_2067 : _GEN_1967; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2093 = _T_202 & oparg_2[5] ? _GEN_2068 : _GEN_1968; // @[NulCtrlMP.scala 557:48]
  wire [63:0] _GEN_2094 = _T_202 & oparg_2[5] ? _GEN_2073 : _GEN_1973; // @[NulCtrlMP.scala 557:48]
  wire [63:0] _GEN_2095 = _T_202 & oparg_2[5] ? _GEN_2074 : _GEN_1974; // @[NulCtrlMP.scala 557:48]
  wire [63:0] _GEN_2096 = _T_202 & oparg_2[5] ? _GEN_2075 : _GEN_1975; // @[NulCtrlMP.scala 557:48]
  wire [63:0] _GEN_2097 = _T_202 & oparg_2[5] ? _GEN_2076 : _GEN_1976; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2098 = _T_202 & oparg_2[5] ? _GEN_2033 : _GEN_1923; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2099 = _T_202 & oparg_2[5] ? _GEN_2034 : _GEN_1924; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2100 = _T_202 & oparg_2[5] ? _GEN_2035 : _GEN_1925; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2101 = _T_202 & oparg_2[5] ? _GEN_2036 : _GEN_1926; // @[NulCtrlMP.scala 557:48]
  wire [31:0] _GEN_2102 = _T_202 & oparg_2[5] ? _GEN_2037 : _GEN_1927; // @[NulCtrlMP.scala 557:48]
  wire [31:0] _GEN_2103 = _T_202 & oparg_2[5] ? _GEN_2038 : _GEN_1928; // @[NulCtrlMP.scala 557:48]
  wire [31:0] _GEN_2104 = _T_202 & oparg_2[5] ? _GEN_2039 : _GEN_1929; // @[NulCtrlMP.scala 557:48]
  wire [31:0] _GEN_2105 = _T_202 & oparg_2[5] ? _GEN_2040 : _GEN_1930; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2106 = _T_202 & oparg_2[5] ? _GEN_2047 : _GEN_1931; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2107 = _T_202 & oparg_2[5] ? _GEN_2048 : _GEN_1932; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2108 = _T_202 & oparg_2[5] ? _GEN_2049 : _GEN_1933; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2109 = _T_202 & oparg_2[5] ? _GEN_2050 : _GEN_1934; // @[NulCtrlMP.scala 557:48]
  wire [4:0] _GEN_2110 = _T_202 & oparg_2[5] ? _GEN_2079 : _GEN_1977; // @[NulCtrlMP.scala 557:48]
  wire  _GEN_2111 = _GEN_145 | _GEN_2080; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2112 = _GEN_146 | _GEN_2081; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2113 = _GEN_147 | _GEN_2082; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2114 = _GEN_148 | _GEN_2083; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_2115 = 2'h0 == opidx ? 5'h5 : _GEN_2084; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2116 = 2'h1 == opidx ? 5'h5 : _GEN_2085; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2117 = 2'h2 == opidx ? 5'h5 : _GEN_2086; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2118 = 2'h3 == opidx ? 5'h5 : _GEN_2087; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_2119 = _T_122 ? _cnt_T : _GEN_2088; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_2120 = _T_122 ? _GEN_1349 : _GEN_2089; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_2121 = cnt[0] ? _GEN_2111 : _GEN_2080; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2122 = cnt[0] ? _GEN_2112 : _GEN_2081; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2123 = cnt[0] ? _GEN_2113 : _GEN_2082; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2124 = cnt[0] ? _GEN_2114 : _GEN_2083; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2125 = cnt[0] ? _GEN_2115 : _GEN_2084; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2126 = cnt[0] ? _GEN_2116 : _GEN_2085; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2127 = cnt[0] ? _GEN_2117 : _GEN_2086; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2128 = cnt[0] ? _GEN_2118 : _GEN_2087; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_2129 = cnt[0] ? _GEN_2119 : _GEN_2088; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_2130 = cnt[0] ? _GEN_2120 : _GEN_2089; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2131 = _GEN_145 | _GEN_2121; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2132 = _GEN_146 | _GEN_2122; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2133 = _GEN_147 | _GEN_2123; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2134 = _GEN_148 | _GEN_2124; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_2135 = 2'h0 == opidx ? 5'h6 : _GEN_2125; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2136 = 2'h1 == opidx ? 5'h6 : _GEN_2126; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2137 = 2'h2 == opidx ? 5'h6 : _GEN_2127; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2138 = 2'h3 == opidx ? 5'h6 : _GEN_2128; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_2139 = _T_122 ? _cnt_T : _GEN_2129; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_2140 = _T_122 ? _GEN_1349 : _GEN_1703; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_2141 = cnt[1] ? _GEN_2131 : _GEN_2121; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2142 = cnt[1] ? _GEN_2132 : _GEN_2122; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2143 = cnt[1] ? _GEN_2133 : _GEN_2123; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2144 = cnt[1] ? _GEN_2134 : _GEN_2124; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2145 = cnt[1] ? _GEN_2135 : _GEN_2125; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2146 = cnt[1] ? _GEN_2136 : _GEN_2126; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2147 = cnt[1] ? _GEN_2137 : _GEN_2127; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2148 = cnt[1] ? _GEN_2138 : _GEN_2128; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_2149 = cnt[1] ? _GEN_2139 : _GEN_2129; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_2150 = cnt[1] ? _GEN_2140 : _GEN_1703; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2151 = _GEN_145 | _GEN_2141; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2152 = _GEN_146 | _GEN_2142; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2153 = _GEN_147 | _GEN_2143; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2154 = _GEN_148 | _GEN_2144; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_2155 = 2'h0 == opidx ? 5'h7 : _GEN_2145; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2156 = 2'h1 == opidx ? 5'h7 : _GEN_2146; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2157 = 2'h2 == opidx ? 5'h7 : _GEN_2147; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2158 = 2'h3 == opidx ? 5'h7 : _GEN_2148; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_2159 = _T_122 ? _cnt_T : _GEN_2149; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_2160 = _T_122 ? _GEN_1349 : regback_2; // @[NulCtrlMP.scala 353:36 355:17 346:26]
  wire  _GEN_2161 = cnt[2] ? _GEN_2151 : _GEN_2141; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2162 = cnt[2] ? _GEN_2152 : _GEN_2142; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2163 = cnt[2] ? _GEN_2153 : _GEN_2143; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2164 = cnt[2] ? _GEN_2154 : _GEN_2144; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2165 = cnt[2] ? _GEN_2155 : _GEN_2145; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2166 = cnt[2] ? _GEN_2156 : _GEN_2146; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2167 = cnt[2] ? _GEN_2157 : _GEN_2147; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2168 = cnt[2] ? _GEN_2158 : _GEN_2148; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_2169 = cnt[2] ? _GEN_2159 : _GEN_2149; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_2170 = cnt[2] ? _GEN_2160 : regback_2; // @[NulCtrlMP.scala 346:26 408:32]
  wire  _GEN_2171 = _GEN_145 | _GEN_2098; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2172 = _GEN_146 | _GEN_2099; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2173 = _GEN_147 | _GEN_2100; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2174 = _GEN_148 | _GEN_2101; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2175 = 2'h0 == opidx ? 32'h342022f3 : _GEN_2102; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2176 = 2'h1 == opidx ? 32'h342022f3 : _GEN_2103; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2177 = 2'h2 == opidx ? 32'h342022f3 : _GEN_2104; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2178 = 2'h3 == opidx ? 32'h342022f3 : _GEN_2105; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2179 = _GEN_1180 ? _cnt_T : _GEN_2169; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2180 = cnt[3] ? _GEN_2171 : _GEN_2098; // @[NulCtrlMP.scala 571:22]
  wire  _GEN_2181 = cnt[3] ? _GEN_2172 : _GEN_2099; // @[NulCtrlMP.scala 571:22]
  wire  _GEN_2182 = cnt[3] ? _GEN_2173 : _GEN_2100; // @[NulCtrlMP.scala 571:22]
  wire  _GEN_2183 = cnt[3] ? _GEN_2174 : _GEN_2101; // @[NulCtrlMP.scala 571:22]
  wire [31:0] _GEN_2184 = cnt[3] ? _GEN_2175 : _GEN_2102; // @[NulCtrlMP.scala 571:22]
  wire [31:0] _GEN_2185 = cnt[3] ? _GEN_2176 : _GEN_2103; // @[NulCtrlMP.scala 571:22]
  wire [31:0] _GEN_2186 = cnt[3] ? _GEN_2177 : _GEN_2104; // @[NulCtrlMP.scala 571:22]
  wire [31:0] _GEN_2187 = cnt[3] ? _GEN_2178 : _GEN_2105; // @[NulCtrlMP.scala 571:22]
  wire [128:0] _GEN_2188 = cnt[3] ? _GEN_2179 : _GEN_2169; // @[NulCtrlMP.scala 571:22]
  wire  _GEN_2189 = _GEN_145 | _GEN_2180; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2190 = _GEN_146 | _GEN_2181; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2191 = _GEN_147 | _GEN_2182; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2192 = _GEN_148 | _GEN_2183; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2193 = 2'h0 == opidx ? 32'h34102373 : _GEN_2184; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2194 = 2'h1 == opidx ? 32'h34102373 : _GEN_2185; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2195 = 2'h2 == opidx ? 32'h34102373 : _GEN_2186; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2196 = 2'h3 == opidx ? 32'h34102373 : _GEN_2187; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2197 = _GEN_1180 ? _cnt_T : _GEN_2188; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2198 = cnt[4] ? _GEN_2189 : _GEN_2180; // @[NulCtrlMP.scala 572:22]
  wire  _GEN_2199 = cnt[4] ? _GEN_2190 : _GEN_2181; // @[NulCtrlMP.scala 572:22]
  wire  _GEN_2200 = cnt[4] ? _GEN_2191 : _GEN_2182; // @[NulCtrlMP.scala 572:22]
  wire  _GEN_2201 = cnt[4] ? _GEN_2192 : _GEN_2183; // @[NulCtrlMP.scala 572:22]
  wire [31:0] _GEN_2202 = cnt[4] ? _GEN_2193 : _GEN_2184; // @[NulCtrlMP.scala 572:22]
  wire [31:0] _GEN_2203 = cnt[4] ? _GEN_2194 : _GEN_2185; // @[NulCtrlMP.scala 572:22]
  wire [31:0] _GEN_2204 = cnt[4] ? _GEN_2195 : _GEN_2186; // @[NulCtrlMP.scala 572:22]
  wire [31:0] _GEN_2205 = cnt[4] ? _GEN_2196 : _GEN_2187; // @[NulCtrlMP.scala 572:22]
  wire [128:0] _GEN_2206 = cnt[4] ? _GEN_2197 : _GEN_2188; // @[NulCtrlMP.scala 572:22]
  wire  _GEN_2207 = _GEN_145 | _GEN_2198; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2208 = _GEN_146 | _GEN_2199; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2209 = _GEN_147 | _GEN_2200; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2210 = _GEN_148 | _GEN_2201; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2211 = 2'h0 == opidx ? 32'h343023f3 : _GEN_2202; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2212 = 2'h1 == opidx ? 32'h343023f3 : _GEN_2203; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2213 = 2'h2 == opidx ? 32'h343023f3 : _GEN_2204; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2214 = 2'h3 == opidx ? 32'h343023f3 : _GEN_2205; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2215 = _GEN_1180 ? _cnt_T : _GEN_2206; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2216 = cnt[5] ? _GEN_2207 : _GEN_2198; // @[NulCtrlMP.scala 573:22]
  wire  _GEN_2217 = cnt[5] ? _GEN_2208 : _GEN_2199; // @[NulCtrlMP.scala 573:22]
  wire  _GEN_2218 = cnt[5] ? _GEN_2209 : _GEN_2200; // @[NulCtrlMP.scala 573:22]
  wire  _GEN_2219 = cnt[5] ? _GEN_2210 : _GEN_2201; // @[NulCtrlMP.scala 573:22]
  wire [31:0] _GEN_2220 = cnt[5] ? _GEN_2211 : _GEN_2202; // @[NulCtrlMP.scala 573:22]
  wire [31:0] _GEN_2221 = cnt[5] ? _GEN_2212 : _GEN_2203; // @[NulCtrlMP.scala 573:22]
  wire [31:0] _GEN_2222 = cnt[5] ? _GEN_2213 : _GEN_2204; // @[NulCtrlMP.scala 573:22]
  wire [31:0] _GEN_2223 = cnt[5] ? _GEN_2214 : _GEN_2205; // @[NulCtrlMP.scala 573:22]
  wire [128:0] _GEN_2224 = cnt[5] ? _GEN_2215 : _GEN_2206; // @[NulCtrlMP.scala 573:22]
  wire  _GEN_2225 = _GEN_145 | _GEN_2106; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_2226 = _GEN_146 | _GEN_2107; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_2227 = _GEN_147 | _GEN_2108; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_2228 = _GEN_148 | _GEN_2109; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_2229 = ~_GEN_1252 ? _cnt_T : _GEN_2224; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_2230 = cnt[6] ? _GEN_2225 : _GEN_2106; // @[NulCtrlMP.scala 574:22]
  wire  _GEN_2231 = cnt[6] ? _GEN_2226 : _GEN_2107; // @[NulCtrlMP.scala 574:22]
  wire  _GEN_2232 = cnt[6] ? _GEN_2227 : _GEN_2108; // @[NulCtrlMP.scala 574:22]
  wire  _GEN_2233 = cnt[6] ? _GEN_2228 : _GEN_2109; // @[NulCtrlMP.scala 574:22]
  wire [128:0] _GEN_2234 = cnt[6] ? _GEN_2229 : _GEN_2224; // @[NulCtrlMP.scala 574:22]
  wire  _GEN_2235 = _GEN_145 | _GEN_2161; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_2236 = _GEN_146 | _GEN_2162; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_2237 = _GEN_147 | _GEN_2163; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_2238 = _GEN_148 | _GEN_2164; // @[NulCtrlMP.scala 359:{27,27}]
  wire [4:0] _GEN_2239 = 2'h0 == opidx ? 5'h5 : _GEN_2165; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_2240 = 2'h1 == opidx ? 5'h5 : _GEN_2166; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_2241 = 2'h2 == opidx ? 5'h5 : _GEN_2167; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_2242 = 2'h3 == opidx ? 5'h5 : _GEN_2168; // @[NulCtrlMP.scala 360:{28,28}]
  wire [128:0] _GEN_2243 = _T_122 ? _cnt_T : _GEN_2234; // @[NulCtrlMP.scala 361:36 362:17]
  wire [7:0] _GEN_2244 = _T_122 ? _GEN_1349[7:0] : _GEN_1796; // @[NulCtrlMP.scala 361:36 364:33]
  wire  _GEN_2245 = cnt[7] ? _GEN_2235 : _GEN_2161; // @[NulCtrlMP.scala 575:22]
  wire  _GEN_2246 = cnt[7] ? _GEN_2236 : _GEN_2162; // @[NulCtrlMP.scala 575:22]
  wire  _GEN_2247 = cnt[7] ? _GEN_2237 : _GEN_2163; // @[NulCtrlMP.scala 575:22]
  wire  _GEN_2248 = cnt[7] ? _GEN_2238 : _GEN_2164; // @[NulCtrlMP.scala 575:22]
  wire [4:0] _GEN_2249 = cnt[7] ? _GEN_2239 : _GEN_2165; // @[NulCtrlMP.scala 575:22]
  wire [4:0] _GEN_2250 = cnt[7] ? _GEN_2240 : _GEN_2166; // @[NulCtrlMP.scala 575:22]
  wire [4:0] _GEN_2251 = cnt[7] ? _GEN_2241 : _GEN_2167; // @[NulCtrlMP.scala 575:22]
  wire [4:0] _GEN_2252 = cnt[7] ? _GEN_2242 : _GEN_2168; // @[NulCtrlMP.scala 575:22]
  wire [128:0] _GEN_2253 = cnt[7] ? _GEN_2243 : _GEN_2234; // @[NulCtrlMP.scala 575:22]
  wire [7:0] _GEN_2254 = cnt[7] ? _GEN_2244 : _GEN_1796; // @[NulCtrlMP.scala 575:22]
  wire  _GEN_2255 = _GEN_145 | _GEN_2245; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_2256 = _GEN_146 | _GEN_2246; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_2257 = _GEN_147 | _GEN_2247; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_2258 = _GEN_148 | _GEN_2248; // @[NulCtrlMP.scala 359:{27,27}]
  wire [4:0] _GEN_2259 = 2'h0 == opidx ? 5'h6 : _GEN_2249; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_2260 = 2'h1 == opidx ? 5'h6 : _GEN_2250; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_2261 = 2'h2 == opidx ? 5'h6 : _GEN_2251; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_2262 = 2'h3 == opidx ? 5'h6 : _GEN_2252; // @[NulCtrlMP.scala 360:{28,28}]
  wire [128:0] _GEN_2263 = _T_122 ? _cnt_T : _GEN_2253; // @[NulCtrlMP.scala 361:36 362:17]
  wire [7:0] _GEN_2264 = _T_122 ? _GEN_1349[7:0] : _GEN_1935; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_2265 = _T_122 ? _GEN_1349[15:8] : _GEN_1936; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_2266 = _T_122 ? _GEN_1349[23:16] : _GEN_1937; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_2267 = _T_122 ? _GEN_1349[31:24] : _GEN_1938; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_2268 = _T_122 ? _GEN_1349[39:32] : _GEN_1939; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_2269 = _T_122 ? _GEN_1349[47:40] : _GEN_1940; // @[NulCtrlMP.scala 361:36 364:33]
  wire  _GEN_2270 = cnt[8] ? _GEN_2255 : _GEN_2245; // @[NulCtrlMP.scala 576:22]
  wire  _GEN_2271 = cnt[8] ? _GEN_2256 : _GEN_2246; // @[NulCtrlMP.scala 576:22]
  wire  _GEN_2272 = cnt[8] ? _GEN_2257 : _GEN_2247; // @[NulCtrlMP.scala 576:22]
  wire  _GEN_2273 = cnt[8] ? _GEN_2258 : _GEN_2248; // @[NulCtrlMP.scala 576:22]
  wire [4:0] _GEN_2274 = cnt[8] ? _GEN_2259 : _GEN_2249; // @[NulCtrlMP.scala 576:22]
  wire [4:0] _GEN_2275 = cnt[8] ? _GEN_2260 : _GEN_2250; // @[NulCtrlMP.scala 576:22]
  wire [4:0] _GEN_2276 = cnt[8] ? _GEN_2261 : _GEN_2251; // @[NulCtrlMP.scala 576:22]
  wire [4:0] _GEN_2277 = cnt[8] ? _GEN_2262 : _GEN_2252; // @[NulCtrlMP.scala 576:22]
  wire [128:0] _GEN_2278 = cnt[8] ? _GEN_2263 : _GEN_2253; // @[NulCtrlMP.scala 576:22]
  wire [7:0] _GEN_2279 = cnt[8] ? _GEN_2264 : _GEN_1935; // @[NulCtrlMP.scala 576:22]
  wire [7:0] _GEN_2280 = cnt[8] ? _GEN_2265 : _GEN_1936; // @[NulCtrlMP.scala 576:22]
  wire [7:0] _GEN_2281 = cnt[8] ? _GEN_2266 : _GEN_1937; // @[NulCtrlMP.scala 576:22]
  wire [7:0] _GEN_2282 = cnt[8] ? _GEN_2267 : _GEN_1938; // @[NulCtrlMP.scala 576:22]
  wire [7:0] _GEN_2283 = cnt[8] ? _GEN_2268 : _GEN_1939; // @[NulCtrlMP.scala 576:22]
  wire [7:0] _GEN_2284 = cnt[8] ? _GEN_2269 : _GEN_1940; // @[NulCtrlMP.scala 576:22]
  wire  _GEN_2285 = _GEN_145 | _GEN_2270; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_2286 = _GEN_146 | _GEN_2271; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_2287 = _GEN_147 | _GEN_2272; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_2288 = _GEN_148 | _GEN_2273; // @[NulCtrlMP.scala 359:{27,27}]
  wire [4:0] _GEN_2289 = 2'h0 == opidx ? 5'h7 : _GEN_2274; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_2290 = 2'h1 == opidx ? 5'h7 : _GEN_2275; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_2291 = 2'h2 == opidx ? 5'h7 : _GEN_2276; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_2292 = 2'h3 == opidx ? 5'h7 : _GEN_2277; // @[NulCtrlMP.scala 360:{28,28}]
  wire [128:0] _GEN_2293 = _T_122 ? _cnt_T : _GEN_2278; // @[NulCtrlMP.scala 361:36 362:17]
  wire [7:0] _GEN_2294 = _T_122 ? _GEN_1349[7:0] : _GEN_1941; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_2295 = _T_122 ? _GEN_1349[15:8] : _GEN_1942; // @[NulCtrlMP.scala 361:36 364:33]
  wire [7:0] _GEN_2296 = _T_122 ? _GEN_1349[23:16] : retarg_10; // @[NulCtrlMP.scala 152:25 361:36 364:33]
  wire [7:0] _GEN_2297 = _T_122 ? _GEN_1349[31:24] : retarg_11; // @[NulCtrlMP.scala 152:25 361:36 364:33]
  wire [7:0] _GEN_2298 = _T_122 ? _GEN_1349[39:32] : retarg_12; // @[NulCtrlMP.scala 152:25 361:36 364:33]
  wire [7:0] _GEN_2299 = _T_122 ? _GEN_1349[47:40] : retarg_13; // @[NulCtrlMP.scala 152:25 361:36 364:33]
  wire  _GEN_2300 = cnt[9] ? _GEN_2285 : _GEN_2270; // @[NulCtrlMP.scala 577:22]
  wire  _GEN_2301 = cnt[9] ? _GEN_2286 : _GEN_2271; // @[NulCtrlMP.scala 577:22]
  wire  _GEN_2302 = cnt[9] ? _GEN_2287 : _GEN_2272; // @[NulCtrlMP.scala 577:22]
  wire  _GEN_2303 = cnt[9] ? _GEN_2288 : _GEN_2273; // @[NulCtrlMP.scala 577:22]
  wire [4:0] _GEN_2304 = cnt[9] ? _GEN_2289 : _GEN_2274; // @[NulCtrlMP.scala 577:22]
  wire [4:0] _GEN_2305 = cnt[9] ? _GEN_2290 : _GEN_2275; // @[NulCtrlMP.scala 577:22]
  wire [4:0] _GEN_2306 = cnt[9] ? _GEN_2291 : _GEN_2276; // @[NulCtrlMP.scala 577:22]
  wire [4:0] _GEN_2307 = cnt[9] ? _GEN_2292 : _GEN_2277; // @[NulCtrlMP.scala 577:22]
  wire [128:0] _GEN_2308 = cnt[9] ? _GEN_2293 : _GEN_2278; // @[NulCtrlMP.scala 577:22]
  wire [7:0] _GEN_2309 = cnt[9] ? _GEN_2294 : _GEN_1941; // @[NulCtrlMP.scala 577:22]
  wire [7:0] _GEN_2310 = cnt[9] ? _GEN_2295 : _GEN_1942; // @[NulCtrlMP.scala 577:22]
  wire [7:0] _GEN_2311 = cnt[9] ? _GEN_2296 : retarg_10; // @[NulCtrlMP.scala 577:22 152:25]
  wire [7:0] _GEN_2312 = cnt[9] ? _GEN_2297 : retarg_11; // @[NulCtrlMP.scala 577:22 152:25]
  wire [7:0] _GEN_2313 = cnt[9] ? _GEN_2298 : retarg_12; // @[NulCtrlMP.scala 577:22 152:25]
  wire [7:0] _GEN_2314 = cnt[9] ? _GEN_2299 : retarg_13; // @[NulCtrlMP.scala 577:22 152:25]
  wire  _GEN_2315 = _GEN_145 | _GEN_2090; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2316 = _GEN_146 | _GEN_2091; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2317 = _GEN_147 | _GEN_2092; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2318 = _GEN_148 | _GEN_2093; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_2319 = 2'h0 == opidx ? 5'h5 : _GEN_2304; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2320 = 2'h1 == opidx ? 5'h5 : _GEN_2305; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2321 = 2'h2 == opidx ? 5'h5 : _GEN_2306; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2322 = 2'h3 == opidx ? 5'h5 : _GEN_2307; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_2323 = 2'h0 == opidx ? regback_0 : _GEN_2094; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2324 = 2'h1 == opidx ? regback_0 : _GEN_2095; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2325 = 2'h2 == opidx ? regback_0 : _GEN_2096; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2326 = 2'h3 == opidx ? regback_0 : _GEN_2097; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_2327 = ~_GEN_1128 ? _cnt_T : _GEN_2308; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_2328 = cnt[10] ? _GEN_2315 : _GEN_2090; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2329 = cnt[10] ? _GEN_2316 : _GEN_2091; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2330 = cnt[10] ? _GEN_2317 : _GEN_2092; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2331 = cnt[10] ? _GEN_2318 : _GEN_2093; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2332 = cnt[10] ? _GEN_2319 : _GEN_2304; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2333 = cnt[10] ? _GEN_2320 : _GEN_2305; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2334 = cnt[10] ? _GEN_2321 : _GEN_2306; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2335 = cnt[10] ? _GEN_2322 : _GEN_2307; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2336 = cnt[10] ? _GEN_2323 : _GEN_2094; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2337 = cnt[10] ? _GEN_2324 : _GEN_2095; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2338 = cnt[10] ? _GEN_2325 : _GEN_2096; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2339 = cnt[10] ? _GEN_2326 : _GEN_2097; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_2340 = cnt[10] ? _GEN_2327 : _GEN_2308; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2341 = _GEN_145 | _GEN_2328; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2342 = _GEN_146 | _GEN_2329; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2343 = _GEN_147 | _GEN_2330; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2344 = _GEN_148 | _GEN_2331; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_2345 = 2'h0 == opidx ? 5'h6 : _GEN_2332; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2346 = 2'h1 == opidx ? 5'h6 : _GEN_2333; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2347 = 2'h2 == opidx ? 5'h6 : _GEN_2334; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2348 = 2'h3 == opidx ? 5'h6 : _GEN_2335; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_2349 = 2'h0 == opidx ? regback_1 : _GEN_2336; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2350 = 2'h1 == opidx ? regback_1 : _GEN_2337; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2351 = 2'h2 == opidx ? regback_1 : _GEN_2338; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2352 = 2'h3 == opidx ? regback_1 : _GEN_2339; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_2353 = ~_GEN_1128 ? _cnt_T : _GEN_2340; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_2354 = cnt[11] ? _GEN_2341 : _GEN_2328; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2355 = cnt[11] ? _GEN_2342 : _GEN_2329; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2356 = cnt[11] ? _GEN_2343 : _GEN_2330; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2357 = cnt[11] ? _GEN_2344 : _GEN_2331; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2358 = cnt[11] ? _GEN_2345 : _GEN_2332; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2359 = cnt[11] ? _GEN_2346 : _GEN_2333; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2360 = cnt[11] ? _GEN_2347 : _GEN_2334; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2361 = cnt[11] ? _GEN_2348 : _GEN_2335; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2362 = cnt[11] ? _GEN_2349 : _GEN_2336; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2363 = cnt[11] ? _GEN_2350 : _GEN_2337; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2364 = cnt[11] ? _GEN_2351 : _GEN_2338; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2365 = cnt[11] ? _GEN_2352 : _GEN_2339; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_2366 = cnt[11] ? _GEN_2353 : _GEN_2340; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2367 = _GEN_145 | _GEN_2354; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2368 = _GEN_146 | _GEN_2355; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2369 = _GEN_147 | _GEN_2356; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_2370 = _GEN_148 | _GEN_2357; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_2371 = 2'h0 == opidx ? 5'h7 : _GEN_2358; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2372 = 2'h1 == opidx ? 5'h7 : _GEN_2359; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2373 = 2'h2 == opidx ? 5'h7 : _GEN_2360; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_2374 = 2'h3 == opidx ? 5'h7 : _GEN_2361; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_2375 = 2'h0 == opidx ? regback_2 : _GEN_2362; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2376 = 2'h1 == opidx ? regback_2 : _GEN_2363; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2377 = 2'h2 == opidx ? regback_2 : _GEN_2364; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_2378 = 2'h3 == opidx ? regback_2 : _GEN_2365; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_2379 = ~_GEN_1128 ? _cnt_T : _GEN_2366; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_2380 = cnt[12] ? _GEN_2367 : _GEN_2354; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2381 = cnt[12] ? _GEN_2368 : _GEN_2355; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2382 = cnt[12] ? _GEN_2369 : _GEN_2356; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2383 = cnt[12] ? _GEN_2370 : _GEN_2357; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2384 = cnt[12] ? _GEN_2371 : _GEN_2358; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2385 = cnt[12] ? _GEN_2372 : _GEN_2359; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2386 = cnt[12] ? _GEN_2373 : _GEN_2360; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_2387 = cnt[12] ? _GEN_2374 : _GEN_2361; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2388 = cnt[12] ? _GEN_2375 : _GEN_2362; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2389 = cnt[12] ? _GEN_2376 : _GEN_2363; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2390 = cnt[12] ? _GEN_2377 : _GEN_2364; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_2391 = cnt[12] ? _GEN_2378 : _GEN_2365; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_2392 = cnt[12] ? _GEN_2379 : _GEN_2366; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_2393 = _GEN_145 | _GEN_2300; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2394 = _GEN_146 | _GEN_2301; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2395 = _GEN_147 | _GEN_2302; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2396 = _GEN_148 | _GEN_2303; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_2397 = 2'h0 == opidx ? 5'h11 : _GEN_2384; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2398 = 2'h1 == opidx ? 5'h11 : _GEN_2385; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2399 = 2'h2 == opidx ? 5'h11 : _GEN_2386; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2400 = 2'h3 == opidx ? 5'h11 : _GEN_2387; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_2401 = _T_122 ? _cnt_T : _GEN_2392; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_2402 = _T_122 ? _GEN_1349 : _GEN_2130; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_2403 = cnt[13] ? _GEN_2393 : _GEN_2300; // @[NulCtrlMP.scala 579:23]
  wire  _GEN_2404 = cnt[13] ? _GEN_2394 : _GEN_2301; // @[NulCtrlMP.scala 579:23]
  wire  _GEN_2405 = cnt[13] ? _GEN_2395 : _GEN_2302; // @[NulCtrlMP.scala 579:23]
  wire  _GEN_2406 = cnt[13] ? _GEN_2396 : _GEN_2303; // @[NulCtrlMP.scala 579:23]
  wire [4:0] _GEN_2407 = cnt[13] ? _GEN_2397 : _GEN_2384; // @[NulCtrlMP.scala 579:23]
  wire [4:0] _GEN_2408 = cnt[13] ? _GEN_2398 : _GEN_2385; // @[NulCtrlMP.scala 579:23]
  wire [4:0] _GEN_2409 = cnt[13] ? _GEN_2399 : _GEN_2386; // @[NulCtrlMP.scala 579:23]
  wire [4:0] _GEN_2410 = cnt[13] ? _GEN_2400 : _GEN_2387; // @[NulCtrlMP.scala 579:23]
  wire [128:0] _GEN_2411 = cnt[13] ? _GEN_2401 : _GEN_2392; // @[NulCtrlMP.scala 579:23]
  wire [63:0] _GEN_2412 = cnt[13] ? _GEN_2402 : _GEN_2130; // @[NulCtrlMP.scala 579:23]
  wire  _T_250 = retarg_1 == 8'h8; // @[NulCtrlMP.scala 582:28]
  wire [4:0] _GEN_2419 = _T_250 & regback_0 == 64'h62 ? 5'h18 : 5'h5; // @[NulCtrlMP.scala 587:76 588:23 590:23]
  wire [128:0] _GEN_2420 = cnt[14] ? 129'h1 : _GEN_2411; // @[NulCtrlMP.scala 580:23 581:17]
  wire [4:0] _GEN_2427 = cnt[14] ? _GEN_2419 : _GEN_2110; // @[NulCtrlMP.scala 580:23]
  wire  _GEN_2428 = state == 5'h9 ? _GEN_2403 : _GEN_2080; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2429 = state == 5'h9 ? _GEN_2404 : _GEN_2081; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2430 = state == 5'h9 ? _GEN_2405 : _GEN_2082; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2431 = state == 5'h9 ? _GEN_2406 : _GEN_2083; // @[NulCtrlMP.scala 569:32]
  wire [4:0] _GEN_2432 = state == 5'h9 ? _GEN_2407 : _GEN_2084; // @[NulCtrlMP.scala 569:32]
  wire [4:0] _GEN_2433 = state == 5'h9 ? _GEN_2408 : _GEN_2085; // @[NulCtrlMP.scala 569:32]
  wire [4:0] _GEN_2434 = state == 5'h9 ? _GEN_2409 : _GEN_2086; // @[NulCtrlMP.scala 569:32]
  wire [4:0] _GEN_2435 = state == 5'h9 ? _GEN_2410 : _GEN_2087; // @[NulCtrlMP.scala 569:32]
  wire [128:0] _GEN_2436 = state == 5'h9 ? _GEN_2420 : _GEN_2088; // @[NulCtrlMP.scala 569:32]
  wire [63:0] _GEN_2437 = state == 5'h9 ? _GEN_2412 : _GEN_2089; // @[NulCtrlMP.scala 569:32]
  wire [63:0] _GEN_2438 = state == 5'h9 ? _GEN_2150 : _GEN_1703; // @[NulCtrlMP.scala 569:32]
  wire [63:0] _GEN_2439 = state == 5'h9 ? _GEN_2170 : regback_2; // @[NulCtrlMP.scala 346:26 569:32]
  wire  _GEN_2440 = state == 5'h9 ? _GEN_2216 : _GEN_2098; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2441 = state == 5'h9 ? _GEN_2217 : _GEN_2099; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2442 = state == 5'h9 ? _GEN_2218 : _GEN_2100; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2443 = state == 5'h9 ? _GEN_2219 : _GEN_2101; // @[NulCtrlMP.scala 569:32]
  wire [31:0] _GEN_2444 = state == 5'h9 ? _GEN_2220 : _GEN_2102; // @[NulCtrlMP.scala 569:32]
  wire [31:0] _GEN_2445 = state == 5'h9 ? _GEN_2221 : _GEN_2103; // @[NulCtrlMP.scala 569:32]
  wire [31:0] _GEN_2446 = state == 5'h9 ? _GEN_2222 : _GEN_2104; // @[NulCtrlMP.scala 569:32]
  wire [31:0] _GEN_2447 = state == 5'h9 ? _GEN_2223 : _GEN_2105; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2448 = state == 5'h9 ? _GEN_2230 : _GEN_2106; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2449 = state == 5'h9 ? _GEN_2231 : _GEN_2107; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2450 = state == 5'h9 ? _GEN_2232 : _GEN_2108; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2451 = state == 5'h9 ? _GEN_2233 : _GEN_2109; // @[NulCtrlMP.scala 569:32]
  wire [7:0] _GEN_2452 = state == 5'h9 ? _GEN_2254 : _GEN_1796; // @[NulCtrlMP.scala 569:32]
  wire [7:0] _GEN_2453 = state == 5'h9 ? _GEN_2279 : _GEN_1935; // @[NulCtrlMP.scala 569:32]
  wire [7:0] _GEN_2454 = state == 5'h9 ? _GEN_2280 : _GEN_1936; // @[NulCtrlMP.scala 569:32]
  wire [7:0] _GEN_2455 = state == 5'h9 ? _GEN_2281 : _GEN_1937; // @[NulCtrlMP.scala 569:32]
  wire [7:0] _GEN_2456 = state == 5'h9 ? _GEN_2282 : _GEN_1938; // @[NulCtrlMP.scala 569:32]
  wire [7:0] _GEN_2457 = state == 5'h9 ? _GEN_2283 : _GEN_1939; // @[NulCtrlMP.scala 569:32]
  wire [7:0] _GEN_2458 = state == 5'h9 ? _GEN_2284 : _GEN_1940; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2465 = state == 5'h9 ? _GEN_2380 : _GEN_2090; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2466 = state == 5'h9 ? _GEN_2381 : _GEN_2091; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2467 = state == 5'h9 ? _GEN_2382 : _GEN_2092; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2468 = state == 5'h9 ? _GEN_2383 : _GEN_2093; // @[NulCtrlMP.scala 569:32]
  wire [63:0] _GEN_2469 = state == 5'h9 ? _GEN_2388 : _GEN_2094; // @[NulCtrlMP.scala 569:32]
  wire [63:0] _GEN_2470 = state == 5'h9 ? _GEN_2389 : _GEN_2095; // @[NulCtrlMP.scala 569:32]
  wire [63:0] _GEN_2471 = state == 5'h9 ? _GEN_2390 : _GEN_2096; // @[NulCtrlMP.scala 569:32]
  wire [63:0] _GEN_2472 = state == 5'h9 ? _GEN_2391 : _GEN_2097; // @[NulCtrlMP.scala 569:32]
  wire [4:0] _GEN_2473 = state == 5'h9 ? _GEN_2427 : _GEN_2110; // @[NulCtrlMP.scala 569:32]
  wire  _GEN_2474 = _GEN_145 | _GEN_2428; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2475 = _GEN_146 | _GEN_2429; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2476 = _GEN_147 | _GEN_2430; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2477 = _GEN_148 | _GEN_2431; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_2478 = 2'h0 == opidx ? 5'ha : _GEN_2432; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2479 = 2'h1 == opidx ? 5'ha : _GEN_2433; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2480 = 2'h2 == opidx ? 5'ha : _GEN_2434; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2481 = 2'h3 == opidx ? 5'ha : _GEN_2435; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_2482 = _T_122 ? _cnt_T : _GEN_2436; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_2483 = _T_122 ? _GEN_1349 : {{16'd0}, hfutex_match_reg}; // @[NulCtrlMP.scala 353:36 355:17 164:35]
  wire  _GEN_2484 = cnt[0] ? _GEN_2474 : _GEN_2428; // @[NulCtrlMP.scala 596:22]
  wire  _GEN_2485 = cnt[0] ? _GEN_2475 : _GEN_2429; // @[NulCtrlMP.scala 596:22]
  wire  _GEN_2486 = cnt[0] ? _GEN_2476 : _GEN_2430; // @[NulCtrlMP.scala 596:22]
  wire  _GEN_2487 = cnt[0] ? _GEN_2477 : _GEN_2431; // @[NulCtrlMP.scala 596:22]
  wire [4:0] _GEN_2488 = cnt[0] ? _GEN_2478 : _GEN_2432; // @[NulCtrlMP.scala 596:22]
  wire [4:0] _GEN_2489 = cnt[0] ? _GEN_2479 : _GEN_2433; // @[NulCtrlMP.scala 596:22]
  wire [4:0] _GEN_2490 = cnt[0] ? _GEN_2480 : _GEN_2434; // @[NulCtrlMP.scala 596:22]
  wire [4:0] _GEN_2491 = cnt[0] ? _GEN_2481 : _GEN_2435; // @[NulCtrlMP.scala 596:22]
  wire [128:0] _GEN_2492 = cnt[0] ? _GEN_2482 : _GEN_2436; // @[NulCtrlMP.scala 596:22]
  wire [63:0] _GEN_2493 = cnt[0] ? _GEN_2483 : {{16'd0}, hfutex_match_reg}; // @[NulCtrlMP.scala 596:22 164:35]
  wire  _GEN_2494 = _GEN_145 | _GEN_2484; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2495 = _GEN_146 | _GEN_2485; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2496 = _GEN_147 | _GEN_2486; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2497 = _GEN_148 | _GEN_2487; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_2498 = 2'h0 == opidx ? 5'hb : _GEN_2488; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2499 = 2'h1 == opidx ? 5'hb : _GEN_2489; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2500 = 2'h2 == opidx ? 5'hb : _GEN_2490; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2501 = 2'h3 == opidx ? 5'hb : _GEN_2491; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_2502 = _T_122 ? _cnt_T : _GEN_2492; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_2503 = _T_122 ? _GEN_1349 : _GEN_2438; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_2504 = cnt[1] ? _GEN_2494 : _GEN_2484; // @[NulCtrlMP.scala 597:22]
  wire  _GEN_2505 = cnt[1] ? _GEN_2495 : _GEN_2485; // @[NulCtrlMP.scala 597:22]
  wire  _GEN_2506 = cnt[1] ? _GEN_2496 : _GEN_2486; // @[NulCtrlMP.scala 597:22]
  wire  _GEN_2507 = cnt[1] ? _GEN_2497 : _GEN_2487; // @[NulCtrlMP.scala 597:22]
  wire [4:0] _GEN_2508 = cnt[1] ? _GEN_2498 : _GEN_2488; // @[NulCtrlMP.scala 597:22]
  wire [4:0] _GEN_2509 = cnt[1] ? _GEN_2499 : _GEN_2489; // @[NulCtrlMP.scala 597:22]
  wire [4:0] _GEN_2510 = cnt[1] ? _GEN_2500 : _GEN_2490; // @[NulCtrlMP.scala 597:22]
  wire [4:0] _GEN_2511 = cnt[1] ? _GEN_2501 : _GEN_2491; // @[NulCtrlMP.scala 597:22]
  wire [128:0] _GEN_2512 = cnt[1] ? _GEN_2502 : _GEN_2492; // @[NulCtrlMP.scala 597:22]
  wire [63:0] _GEN_2513 = cnt[1] ? _GEN_2503 : _GEN_2438; // @[NulCtrlMP.scala 597:22]
  wire [128:0] _GEN_2514 = regback_1[6:0] == 7'h1 & hfutex_match_reg != 48'h0 & hfutex_hit ? _cnt_T : 129'h1; // @[NulCtrlMP.scala 599:88 600:21 602:21]
  wire [4:0] _GEN_2515 = regback_1[6:0] == 7'h1 & hfutex_match_reg != 48'h0 & hfutex_hit ? _GEN_2473 : 5'h5; // @[NulCtrlMP.scala 599:88 603:23]
  wire [128:0] _GEN_2516 = cnt[2] ? _GEN_2514 : _GEN_2512; // @[NulCtrlMP.scala 598:22]
  wire [4:0] _GEN_2517 = cnt[2] ? _GEN_2515 : _GEN_2473; // @[NulCtrlMP.scala 598:22]
  wire  _GEN_2518 = _GEN_145 | _GEN_2440; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2519 = _GEN_146 | _GEN_2441; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2520 = _GEN_147 | _GEN_2442; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2521 = _GEN_148 | _GEN_2443; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2522 = 2'h0 == opidx ? 32'h34102573 : _GEN_2444; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2523 = 2'h1 == opidx ? 32'h34102573 : _GEN_2445; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2524 = 2'h2 == opidx ? 32'h34102573 : _GEN_2446; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2525 = 2'h3 == opidx ? 32'h34102573 : _GEN_2447; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2526 = _GEN_1180 ? _cnt_T : _GEN_2516; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2527 = cnt[3] ? _GEN_2518 : _GEN_2440; // @[NulCtrlMP.scala 606:22]
  wire  _GEN_2528 = cnt[3] ? _GEN_2519 : _GEN_2441; // @[NulCtrlMP.scala 606:22]
  wire  _GEN_2529 = cnt[3] ? _GEN_2520 : _GEN_2442; // @[NulCtrlMP.scala 606:22]
  wire  _GEN_2530 = cnt[3] ? _GEN_2521 : _GEN_2443; // @[NulCtrlMP.scala 606:22]
  wire [31:0] _GEN_2531 = cnt[3] ? _GEN_2522 : _GEN_2444; // @[NulCtrlMP.scala 606:22]
  wire [31:0] _GEN_2532 = cnt[3] ? _GEN_2523 : _GEN_2445; // @[NulCtrlMP.scala 606:22]
  wire [31:0] _GEN_2533 = cnt[3] ? _GEN_2524 : _GEN_2446; // @[NulCtrlMP.scala 606:22]
  wire [31:0] _GEN_2534 = cnt[3] ? _GEN_2525 : _GEN_2447; // @[NulCtrlMP.scala 606:22]
  wire [128:0] _GEN_2535 = cnt[3] ? _GEN_2526 : _GEN_2516; // @[NulCtrlMP.scala 606:22]
  wire  _GEN_2536 = _GEN_145 | _GEN_2527; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2537 = _GEN_146 | _GEN_2528; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2538 = _GEN_147 | _GEN_2529; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2539 = _GEN_148 | _GEN_2530; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2540 = 2'h0 == opidx ? 32'h450513 : _GEN_2531; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2541 = 2'h1 == opidx ? 32'h450513 : _GEN_2532; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2542 = 2'h2 == opidx ? 32'h450513 : _GEN_2533; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2543 = 2'h3 == opidx ? 32'h450513 : _GEN_2534; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2544 = _GEN_1180 ? _cnt_T : _GEN_2535; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2545 = cnt[4] ? _GEN_2536 : _GEN_2527; // @[NulCtrlMP.scala 607:22]
  wire  _GEN_2546 = cnt[4] ? _GEN_2537 : _GEN_2528; // @[NulCtrlMP.scala 607:22]
  wire  _GEN_2547 = cnt[4] ? _GEN_2538 : _GEN_2529; // @[NulCtrlMP.scala 607:22]
  wire  _GEN_2548 = cnt[4] ? _GEN_2539 : _GEN_2530; // @[NulCtrlMP.scala 607:22]
  wire [31:0] _GEN_2549 = cnt[4] ? _GEN_2540 : _GEN_2531; // @[NulCtrlMP.scala 607:22]
  wire [31:0] _GEN_2550 = cnt[4] ? _GEN_2541 : _GEN_2532; // @[NulCtrlMP.scala 607:22]
  wire [31:0] _GEN_2551 = cnt[4] ? _GEN_2542 : _GEN_2533; // @[NulCtrlMP.scala 607:22]
  wire [31:0] _GEN_2552 = cnt[4] ? _GEN_2543 : _GEN_2534; // @[NulCtrlMP.scala 607:22]
  wire [128:0] _GEN_2553 = cnt[4] ? _GEN_2544 : _GEN_2535; // @[NulCtrlMP.scala 607:22]
  wire  _GEN_2554 = _GEN_145 | _GEN_2545; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2555 = _GEN_146 | _GEN_2546; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2556 = _GEN_147 | _GEN_2547; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2557 = _GEN_148 | _GEN_2548; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2558 = 2'h0 == opidx ? 32'h34151073 : _GEN_2549; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2559 = 2'h1 == opidx ? 32'h34151073 : _GEN_2550; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2560 = 2'h2 == opidx ? 32'h34151073 : _GEN_2551; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2561 = 2'h3 == opidx ? 32'h34151073 : _GEN_2552; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2562 = _GEN_1180 ? _cnt_T : _GEN_2553; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2563 = cnt[5] ? _GEN_2554 : _GEN_2545; // @[NulCtrlMP.scala 608:22]
  wire  _GEN_2564 = cnt[5] ? _GEN_2555 : _GEN_2546; // @[NulCtrlMP.scala 608:22]
  wire  _GEN_2565 = cnt[5] ? _GEN_2556 : _GEN_2547; // @[NulCtrlMP.scala 608:22]
  wire  _GEN_2566 = cnt[5] ? _GEN_2557 : _GEN_2548; // @[NulCtrlMP.scala 608:22]
  wire [31:0] _GEN_2567 = cnt[5] ? _GEN_2558 : _GEN_2549; // @[NulCtrlMP.scala 608:22]
  wire [31:0] _GEN_2568 = cnt[5] ? _GEN_2559 : _GEN_2550; // @[NulCtrlMP.scala 608:22]
  wire [31:0] _GEN_2569 = cnt[5] ? _GEN_2560 : _GEN_2551; // @[NulCtrlMP.scala 608:22]
  wire [31:0] _GEN_2570 = cnt[5] ? _GEN_2561 : _GEN_2552; // @[NulCtrlMP.scala 608:22]
  wire [128:0] _GEN_2571 = cnt[5] ? _GEN_2562 : _GEN_2553; // @[NulCtrlMP.scala 608:22]
  wire  _GEN_2572 = _GEN_145 | _GEN_2563; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2573 = _GEN_146 | _GEN_2564; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2574 = _GEN_147 | _GEN_2565; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2575 = _GEN_148 | _GEN_2566; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2576 = 2'h0 == opidx ? 32'h300513 : _GEN_2567; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2577 = 2'h1 == opidx ? 32'h300513 : _GEN_2568; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2578 = 2'h2 == opidx ? 32'h300513 : _GEN_2569; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2579 = 2'h3 == opidx ? 32'h300513 : _GEN_2570; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2580 = _GEN_1180 ? _cnt_T : _GEN_2571; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2581 = cnt[6] ? _GEN_2572 : _GEN_2563; // @[NulCtrlMP.scala 609:22]
  wire  _GEN_2582 = cnt[6] ? _GEN_2573 : _GEN_2564; // @[NulCtrlMP.scala 609:22]
  wire  _GEN_2583 = cnt[6] ? _GEN_2574 : _GEN_2565; // @[NulCtrlMP.scala 609:22]
  wire  _GEN_2584 = cnt[6] ? _GEN_2575 : _GEN_2566; // @[NulCtrlMP.scala 609:22]
  wire [31:0] _GEN_2585 = cnt[6] ? _GEN_2576 : _GEN_2567; // @[NulCtrlMP.scala 609:22]
  wire [31:0] _GEN_2586 = cnt[6] ? _GEN_2577 : _GEN_2568; // @[NulCtrlMP.scala 609:22]
  wire [31:0] _GEN_2587 = cnt[6] ? _GEN_2578 : _GEN_2569; // @[NulCtrlMP.scala 609:22]
  wire [31:0] _GEN_2588 = cnt[6] ? _GEN_2579 : _GEN_2570; // @[NulCtrlMP.scala 609:22]
  wire [128:0] _GEN_2589 = cnt[6] ? _GEN_2580 : _GEN_2571; // @[NulCtrlMP.scala 609:22]
  wire  _GEN_2590 = _GEN_145 | _GEN_2581; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2591 = _GEN_146 | _GEN_2582; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2592 = _GEN_147 | _GEN_2583; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2593 = _GEN_148 | _GEN_2584; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2594 = 2'h0 == opidx ? 32'hb51513 : _GEN_2585; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2595 = 2'h1 == opidx ? 32'hb51513 : _GEN_2586; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2596 = 2'h2 == opidx ? 32'hb51513 : _GEN_2587; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2597 = 2'h3 == opidx ? 32'hb51513 : _GEN_2588; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2598 = _GEN_1180 ? _cnt_T : _GEN_2589; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2599 = cnt[7] ? _GEN_2590 : _GEN_2581; // @[NulCtrlMP.scala 610:22]
  wire  _GEN_2600 = cnt[7] ? _GEN_2591 : _GEN_2582; // @[NulCtrlMP.scala 610:22]
  wire  _GEN_2601 = cnt[7] ? _GEN_2592 : _GEN_2583; // @[NulCtrlMP.scala 610:22]
  wire  _GEN_2602 = cnt[7] ? _GEN_2593 : _GEN_2584; // @[NulCtrlMP.scala 610:22]
  wire [31:0] _GEN_2603 = cnt[7] ? _GEN_2594 : _GEN_2585; // @[NulCtrlMP.scala 610:22]
  wire [31:0] _GEN_2604 = cnt[7] ? _GEN_2595 : _GEN_2586; // @[NulCtrlMP.scala 610:22]
  wire [31:0] _GEN_2605 = cnt[7] ? _GEN_2596 : _GEN_2587; // @[NulCtrlMP.scala 610:22]
  wire [31:0] _GEN_2606 = cnt[7] ? _GEN_2597 : _GEN_2588; // @[NulCtrlMP.scala 610:22]
  wire [128:0] _GEN_2607 = cnt[7] ? _GEN_2598 : _GEN_2589; // @[NulCtrlMP.scala 610:22]
  wire  _GEN_2608 = _GEN_145 | _GEN_2599; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2609 = _GEN_146 | _GEN_2600; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2610 = _GEN_147 | _GEN_2601; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2611 = _GEN_148 | _GEN_2602; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2612 = 2'h0 == opidx ? 32'h30053073 : _GEN_2603; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2613 = 2'h1 == opidx ? 32'h30053073 : _GEN_2604; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2614 = 2'h2 == opidx ? 32'h30053073 : _GEN_2605; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2615 = 2'h3 == opidx ? 32'h30053073 : _GEN_2606; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2616 = _GEN_1180 ? _cnt_T : _GEN_2607; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2617 = cnt[8] ? _GEN_2608 : _GEN_2599; // @[NulCtrlMP.scala 611:22]
  wire  _GEN_2618 = cnt[8] ? _GEN_2609 : _GEN_2600; // @[NulCtrlMP.scala 611:22]
  wire  _GEN_2619 = cnt[8] ? _GEN_2610 : _GEN_2601; // @[NulCtrlMP.scala 611:22]
  wire  _GEN_2620 = cnt[8] ? _GEN_2611 : _GEN_2602; // @[NulCtrlMP.scala 611:22]
  wire [31:0] _GEN_2621 = cnt[8] ? _GEN_2612 : _GEN_2603; // @[NulCtrlMP.scala 611:22]
  wire [31:0] _GEN_2622 = cnt[8] ? _GEN_2613 : _GEN_2604; // @[NulCtrlMP.scala 611:22]
  wire [31:0] _GEN_2623 = cnt[8] ? _GEN_2614 : _GEN_2605; // @[NulCtrlMP.scala 611:22]
  wire [31:0] _GEN_2624 = cnt[8] ? _GEN_2615 : _GEN_2606; // @[NulCtrlMP.scala 611:22]
  wire [128:0] _GEN_2625 = cnt[8] ? _GEN_2616 : _GEN_2607; // @[NulCtrlMP.scala 611:22]
  wire  _GEN_2626 = _GEN_145 | _GEN_2617; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2627 = _GEN_146 | _GEN_2618; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2628 = _GEN_147 | _GEN_2619; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2629 = _GEN_148 | _GEN_2620; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2630 = 2'h0 == opidx ? 32'h2537 : _GEN_2621; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2631 = 2'h1 == opidx ? 32'h2537 : _GEN_2622; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2632 = 2'h2 == opidx ? 32'h2537 : _GEN_2623; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2633 = 2'h3 == opidx ? 32'h2537 : _GEN_2624; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2634 = _GEN_1180 ? _cnt_T : _GEN_2625; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2635 = cnt[9] ? _GEN_2626 : _GEN_2617; // @[NulCtrlMP.scala 612:22]
  wire  _GEN_2636 = cnt[9] ? _GEN_2627 : _GEN_2618; // @[NulCtrlMP.scala 612:22]
  wire  _GEN_2637 = cnt[9] ? _GEN_2628 : _GEN_2619; // @[NulCtrlMP.scala 612:22]
  wire  _GEN_2638 = cnt[9] ? _GEN_2629 : _GEN_2620; // @[NulCtrlMP.scala 612:22]
  wire [31:0] _GEN_2639 = cnt[9] ? _GEN_2630 : _GEN_2621; // @[NulCtrlMP.scala 612:22]
  wire [31:0] _GEN_2640 = cnt[9] ? _GEN_2631 : _GEN_2622; // @[NulCtrlMP.scala 612:22]
  wire [31:0] _GEN_2641 = cnt[9] ? _GEN_2632 : _GEN_2623; // @[NulCtrlMP.scala 612:22]
  wire [31:0] _GEN_2642 = cnt[9] ? _GEN_2633 : _GEN_2624; // @[NulCtrlMP.scala 612:22]
  wire [128:0] _GEN_2643 = cnt[9] ? _GEN_2634 : _GEN_2625; // @[NulCtrlMP.scala 612:22]
  wire  _GEN_2644 = _GEN_145 | _GEN_2635; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2645 = _GEN_146 | _GEN_2636; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2646 = _GEN_147 | _GEN_2637; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2647 = _GEN_148 | _GEN_2638; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2648 = 2'h0 == opidx ? 32'h30052073 : _GEN_2639; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2649 = 2'h1 == opidx ? 32'h30052073 : _GEN_2640; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2650 = 2'h2 == opidx ? 32'h30052073 : _GEN_2641; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2651 = 2'h3 == opidx ? 32'h30052073 : _GEN_2642; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2652 = _GEN_1180 ? _cnt_T : _GEN_2643; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2653 = cnt[10] ? _GEN_2644 : _GEN_2635; // @[NulCtrlMP.scala 619:23]
  wire  _GEN_2654 = cnt[10] ? _GEN_2645 : _GEN_2636; // @[NulCtrlMP.scala 619:23]
  wire  _GEN_2655 = cnt[10] ? _GEN_2646 : _GEN_2637; // @[NulCtrlMP.scala 619:23]
  wire  _GEN_2656 = cnt[10] ? _GEN_2647 : _GEN_2638; // @[NulCtrlMP.scala 619:23]
  wire [31:0] _GEN_2657 = cnt[10] ? _GEN_2648 : _GEN_2639; // @[NulCtrlMP.scala 619:23]
  wire [31:0] _GEN_2658 = cnt[10] ? _GEN_2649 : _GEN_2640; // @[NulCtrlMP.scala 619:23]
  wire [31:0] _GEN_2659 = cnt[10] ? _GEN_2650 : _GEN_2641; // @[NulCtrlMP.scala 619:23]
  wire [31:0] _GEN_2660 = cnt[10] ? _GEN_2651 : _GEN_2642; // @[NulCtrlMP.scala 619:23]
  wire [128:0] _GEN_2661 = cnt[10] ? _GEN_2652 : _GEN_2643; // @[NulCtrlMP.scala 619:23]
  wire  _GEN_2662 = _GEN_145 | _GEN_2653; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2663 = _GEN_146 | _GEN_2654; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2664 = _GEN_147 | _GEN_2655; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2665 = _GEN_148 | _GEN_2656; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2666 = 2'h0 == opidx ? 32'h301073 : _GEN_2657; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2667 = 2'h1 == opidx ? 32'h301073 : _GEN_2658; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2668 = 2'h2 == opidx ? 32'h301073 : _GEN_2659; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2669 = 2'h3 == opidx ? 32'h301073 : _GEN_2660; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2670 = _GEN_1180 ? _cnt_T : _GEN_2661; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2671 = cnt[11] ? _GEN_2662 : _GEN_2653; // @[NulCtrlMP.scala 626:23]
  wire  _GEN_2672 = cnt[11] ? _GEN_2663 : _GEN_2654; // @[NulCtrlMP.scala 626:23]
  wire  _GEN_2673 = cnt[11] ? _GEN_2664 : _GEN_2655; // @[NulCtrlMP.scala 626:23]
  wire  _GEN_2674 = cnt[11] ? _GEN_2665 : _GEN_2656; // @[NulCtrlMP.scala 626:23]
  wire [31:0] _GEN_2675 = cnt[11] ? _GEN_2666 : _GEN_2657; // @[NulCtrlMP.scala 626:23]
  wire [31:0] _GEN_2676 = cnt[11] ? _GEN_2667 : _GEN_2658; // @[NulCtrlMP.scala 626:23]
  wire [31:0] _GEN_2677 = cnt[11] ? _GEN_2668 : _GEN_2659; // @[NulCtrlMP.scala 626:23]
  wire [31:0] _GEN_2678 = cnt[11] ? _GEN_2669 : _GEN_2660; // @[NulCtrlMP.scala 626:23]
  wire [128:0] _GEN_2679 = cnt[11] ? _GEN_2670 : _GEN_2661; // @[NulCtrlMP.scala 626:23]
  wire  _GEN_2680 = _GEN_145 | _GEN_2671; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2681 = _GEN_146 | _GEN_2672; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2682 = _GEN_147 | _GEN_2673; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2683 = _GEN_148 | _GEN_2674; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2684 = 2'h0 == opidx ? 32'h330000f : _GEN_2675; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2685 = 2'h1 == opidx ? 32'h330000f : _GEN_2676; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2686 = 2'h2 == opidx ? 32'h330000f : _GEN_2677; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2687 = 2'h3 == opidx ? 32'h330000f : _GEN_2678; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2688 = _GEN_1180 ? _cnt_T : _GEN_2679; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2689 = cnt[12] ? _GEN_2680 : _GEN_2671; // @[NulCtrlMP.scala 633:23]
  wire  _GEN_2690 = cnt[12] ? _GEN_2681 : _GEN_2672; // @[NulCtrlMP.scala 633:23]
  wire  _GEN_2691 = cnt[12] ? _GEN_2682 : _GEN_2673; // @[NulCtrlMP.scala 633:23]
  wire  _GEN_2692 = cnt[12] ? _GEN_2683 : _GEN_2674; // @[NulCtrlMP.scala 633:23]
  wire [31:0] _GEN_2693 = cnt[12] ? _GEN_2684 : _GEN_2675; // @[NulCtrlMP.scala 633:23]
  wire [31:0] _GEN_2694 = cnt[12] ? _GEN_2685 : _GEN_2676; // @[NulCtrlMP.scala 633:23]
  wire [31:0] _GEN_2695 = cnt[12] ? _GEN_2686 : _GEN_2677; // @[NulCtrlMP.scala 633:23]
  wire [31:0] _GEN_2696 = cnt[12] ? _GEN_2687 : _GEN_2678; // @[NulCtrlMP.scala 633:23]
  wire [128:0] _GEN_2697 = cnt[12] ? _GEN_2688 : _GEN_2679; // @[NulCtrlMP.scala 633:23]
  wire  _GEN_2698 = _GEN_145 | _GEN_2689; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2699 = _GEN_146 | _GEN_2690; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2700 = _GEN_147 | _GEN_2691; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2701 = _GEN_148 | _GEN_2692; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2702 = 2'h0 == opidx ? 32'h537 : _GEN_2693; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2703 = 2'h1 == opidx ? 32'h537 : _GEN_2694; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2704 = 2'h2 == opidx ? 32'h537 : _GEN_2695; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2705 = 2'h3 == opidx ? 32'h537 : _GEN_2696; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2706 = _GEN_1180 ? _cnt_T : _GEN_2697; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2707 = cnt[13] ? _GEN_2698 : _GEN_2689; // @[NulCtrlMP.scala 634:23]
  wire  _GEN_2708 = cnt[13] ? _GEN_2699 : _GEN_2690; // @[NulCtrlMP.scala 634:23]
  wire  _GEN_2709 = cnt[13] ? _GEN_2700 : _GEN_2691; // @[NulCtrlMP.scala 634:23]
  wire  _GEN_2710 = cnt[13] ? _GEN_2701 : _GEN_2692; // @[NulCtrlMP.scala 634:23]
  wire [31:0] _GEN_2711 = cnt[13] ? _GEN_2702 : _GEN_2693; // @[NulCtrlMP.scala 634:23]
  wire [31:0] _GEN_2712 = cnt[13] ? _GEN_2703 : _GEN_2694; // @[NulCtrlMP.scala 634:23]
  wire [31:0] _GEN_2713 = cnt[13] ? _GEN_2704 : _GEN_2695; // @[NulCtrlMP.scala 634:23]
  wire [31:0] _GEN_2714 = cnt[13] ? _GEN_2705 : _GEN_2696; // @[NulCtrlMP.scala 634:23]
  wire [128:0] _GEN_2715 = cnt[13] ? _GEN_2706 : _GEN_2697; // @[NulCtrlMP.scala 634:23]
  wire  _GEN_2716 = _GEN_145 | _GEN_2448; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_2717 = _GEN_146 | _GEN_2449; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_2718 = _GEN_147 | _GEN_2450; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_2719 = _GEN_148 | _GEN_2451; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_2720 = ~_GEN_1252 ? _cnt_T : _GEN_2715; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_2721 = cnt[14] ? _GEN_2716 : _GEN_2448; // @[NulCtrlMP.scala 635:23]
  wire  _GEN_2722 = cnt[14] ? _GEN_2717 : _GEN_2449; // @[NulCtrlMP.scala 635:23]
  wire  _GEN_2723 = cnt[14] ? _GEN_2718 : _GEN_2450; // @[NulCtrlMP.scala 635:23]
  wire  _GEN_2724 = cnt[14] ? _GEN_2719 : _GEN_2451; // @[NulCtrlMP.scala 635:23]
  wire [128:0] _GEN_2725 = cnt[14] ? _GEN_2720 : _GEN_2715; // @[NulCtrlMP.scala 635:23]
  wire  _GEN_2730 = _GEN_145 | _GEN_2707; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2731 = _GEN_146 | _GEN_2708; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2732 = _GEN_147 | _GEN_2709; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2733 = _GEN_148 | _GEN_2710; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2734 = 2'h0 == opidx ? 32'h30200073 : _GEN_2711; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2735 = 2'h1 == opidx ? 32'h30200073 : _GEN_2712; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2736 = 2'h2 == opidx ? 32'h30200073 : _GEN_2713; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2737 = 2'h3 == opidx ? 32'h30200073 : _GEN_2714; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2738 = _GEN_1180 ? _cnt_T : _GEN_2725; // @[NulCtrlMP.scala 396:36 397:17]
  wire [1:0] _GEN_2739 = 2'h0 == opidx ? 2'h3 : _GEN_1020; // @[NulCtrlMP.scala 640:{34,34}]
  wire [1:0] _GEN_2740 = 2'h1 == opidx ? 2'h3 : _GEN_1021; // @[NulCtrlMP.scala 640:{34,34}]
  wire [1:0] _GEN_2741 = 2'h2 == opidx ? 2'h3 : _GEN_1022; // @[NulCtrlMP.scala 640:{34,34}]
  wire [1:0] _GEN_2742 = 2'h3 == opidx ? 2'h3 : _GEN_1023; // @[NulCtrlMP.scala 640:{34,34}]
  wire [1:0] _GEN_2743 = _GEN_1180 ? _GEN_2739 : _GEN_1020; // @[NulCtrlMP.scala 639:40]
  wire [1:0] _GEN_2744 = _GEN_1180 ? _GEN_2740 : _GEN_1021; // @[NulCtrlMP.scala 639:40]
  wire [1:0] _GEN_2745 = _GEN_1180 ? _GEN_2741 : _GEN_1022; // @[NulCtrlMP.scala 639:40]
  wire [1:0] _GEN_2746 = _GEN_1180 ? _GEN_2742 : _GEN_1023; // @[NulCtrlMP.scala 639:40]
  wire  _GEN_2747 = cnt[15] & _GEN_145; // @[NulCtrlMP.scala 636:23 51:33]
  wire  _GEN_2748 = cnt[15] & _GEN_146; // @[NulCtrlMP.scala 636:23 51:33]
  wire  _GEN_2749 = cnt[15] & _GEN_147; // @[NulCtrlMP.scala 636:23 51:33]
  wire  _GEN_2750 = cnt[15] & _GEN_148; // @[NulCtrlMP.scala 636:23 51:33]
  wire  _GEN_2751 = cnt[15] ? _GEN_2730 : _GEN_2707; // @[NulCtrlMP.scala 636:23]
  wire  _GEN_2752 = cnt[15] ? _GEN_2731 : _GEN_2708; // @[NulCtrlMP.scala 636:23]
  wire  _GEN_2753 = cnt[15] ? _GEN_2732 : _GEN_2709; // @[NulCtrlMP.scala 636:23]
  wire  _GEN_2754 = cnt[15] ? _GEN_2733 : _GEN_2710; // @[NulCtrlMP.scala 636:23]
  wire [31:0] _GEN_2755 = cnt[15] ? _GEN_2734 : _GEN_2711; // @[NulCtrlMP.scala 636:23]
  wire [31:0] _GEN_2756 = cnt[15] ? _GEN_2735 : _GEN_2712; // @[NulCtrlMP.scala 636:23]
  wire [31:0] _GEN_2757 = cnt[15] ? _GEN_2736 : _GEN_2713; // @[NulCtrlMP.scala 636:23]
  wire [31:0] _GEN_2758 = cnt[15] ? _GEN_2737 : _GEN_2714; // @[NulCtrlMP.scala 636:23]
  wire [128:0] _GEN_2759 = cnt[15] ? _GEN_2738 : _GEN_2725; // @[NulCtrlMP.scala 636:23]
  wire [1:0] _GEN_2760 = cnt[15] ? _GEN_2743 : _GEN_1020; // @[NulCtrlMP.scala 636:23]
  wire [1:0] _GEN_2761 = cnt[15] ? _GEN_2744 : _GEN_1021; // @[NulCtrlMP.scala 636:23]
  wire [1:0] _GEN_2762 = cnt[15] ? _GEN_2745 : _GEN_1022; // @[NulCtrlMP.scala 636:23]
  wire [1:0] _GEN_2763 = cnt[15] ? _GEN_2746 : _GEN_1023; // @[NulCtrlMP.scala 636:23]
  wire  _GEN_2764 = _GEN_145 | _GEN_2721; // @[NulCtrlMP.scala 644:{34,34}]
  wire  _GEN_2765 = _GEN_146 | _GEN_2722; // @[NulCtrlMP.scala 644:{34,34}]
  wire  _GEN_2766 = _GEN_147 | _GEN_2723; // @[NulCtrlMP.scala 644:{34,34}]
  wire  _GEN_2767 = _GEN_148 | _GEN_2724; // @[NulCtrlMP.scala 644:{34,34}]
  wire  _GEN_2768 = cnt[16] ? _GEN_2764 : _GEN_2721; // @[NulCtrlMP.scala 643:23]
  wire  _GEN_2769 = cnt[16] ? _GEN_2765 : _GEN_2722; // @[NulCtrlMP.scala 643:23]
  wire  _GEN_2770 = cnt[16] ? _GEN_2766 : _GEN_2723; // @[NulCtrlMP.scala 643:23]
  wire  _GEN_2771 = cnt[16] ? _GEN_2767 : _GEN_2724; // @[NulCtrlMP.scala 643:23]
  wire [128:0] _GEN_2772 = cnt[16] ? _cnt_T : _GEN_2759; // @[NulCtrlMP.scala 643:23 645:17]
  wire [128:0] _GEN_2773 = cnt[17] ? 129'h1 : _GEN_2772; // @[NulCtrlMP.scala 647:23 648:17]
  wire [4:0] _GEN_2774 = cnt[17] ? 5'h8 : _GEN_2517; // @[NulCtrlMP.scala 647:23 649:19]
  wire  _GEN_2775 = state == 5'h18 ? _GEN_2504 : _GEN_2428; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2776 = state == 5'h18 ? _GEN_2505 : _GEN_2429; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2777 = state == 5'h18 ? _GEN_2506 : _GEN_2430; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2778 = state == 5'h18 ? _GEN_2507 : _GEN_2431; // @[NulCtrlMP.scala 595:34]
  wire [4:0] _GEN_2779 = state == 5'h18 ? _GEN_2508 : _GEN_2432; // @[NulCtrlMP.scala 595:34]
  wire [4:0] _GEN_2780 = state == 5'h18 ? _GEN_2509 : _GEN_2433; // @[NulCtrlMP.scala 595:34]
  wire [4:0] _GEN_2781 = state == 5'h18 ? _GEN_2510 : _GEN_2434; // @[NulCtrlMP.scala 595:34]
  wire [4:0] _GEN_2782 = state == 5'h18 ? _GEN_2511 : _GEN_2435; // @[NulCtrlMP.scala 595:34]
  wire [128:0] _GEN_2783 = state == 5'h18 ? _GEN_2773 : _GEN_2436; // @[NulCtrlMP.scala 595:34]
  wire [63:0] _GEN_2784 = state == 5'h18 ? _GEN_2493 : {{16'd0}, hfutex_match_reg}; // @[NulCtrlMP.scala 595:34 164:35]
  wire [63:0] _GEN_2785 = state == 5'h18 ? _GEN_2513 : _GEN_2438; // @[NulCtrlMP.scala 595:34]
  wire [4:0] _GEN_2786 = state == 5'h18 ? _GEN_2774 : _GEN_2473; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2787 = state == 5'h18 ? _GEN_2751 : _GEN_2440; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2788 = state == 5'h18 ? _GEN_2752 : _GEN_2441; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2789 = state == 5'h18 ? _GEN_2753 : _GEN_2442; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2790 = state == 5'h18 ? _GEN_2754 : _GEN_2443; // @[NulCtrlMP.scala 595:34]
  wire [31:0] _GEN_2791 = state == 5'h18 ? _GEN_2755 : _GEN_2444; // @[NulCtrlMP.scala 595:34]
  wire [31:0] _GEN_2792 = state == 5'h18 ? _GEN_2756 : _GEN_2445; // @[NulCtrlMP.scala 595:34]
  wire [31:0] _GEN_2793 = state == 5'h18 ? _GEN_2757 : _GEN_2446; // @[NulCtrlMP.scala 595:34]
  wire [31:0] _GEN_2794 = state == 5'h18 ? _GEN_2758 : _GEN_2447; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2795 = state == 5'h18 ? _GEN_2768 : _GEN_2448; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2796 = state == 5'h18 ? _GEN_2769 : _GEN_2449; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2797 = state == 5'h18 ? _GEN_2770 : _GEN_2450; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2798 = state == 5'h18 ? _GEN_2771 : _GEN_2451; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2799 = state == 5'h18 & _GEN_2747; // @[NulCtrlMP.scala 51:33 595:34]
  wire  _GEN_2800 = state == 5'h18 & _GEN_2748; // @[NulCtrlMP.scala 51:33 595:34]
  wire  _GEN_2801 = state == 5'h18 & _GEN_2749; // @[NulCtrlMP.scala 51:33 595:34]
  wire  _GEN_2802 = state == 5'h18 & _GEN_2750; // @[NulCtrlMP.scala 51:33 595:34]
  wire [1:0] _GEN_2803 = state == 5'h18 ? _GEN_2760 : _GEN_1020; // @[NulCtrlMP.scala 595:34]
  wire [1:0] _GEN_2804 = state == 5'h18 ? _GEN_2761 : _GEN_1021; // @[NulCtrlMP.scala 595:34]
  wire [1:0] _GEN_2805 = state == 5'h18 ? _GEN_2762 : _GEN_1022; // @[NulCtrlMP.scala 595:34]
  wire [1:0] _GEN_2806 = state == 5'h18 ? _GEN_2763 : _GEN_1023; // @[NulCtrlMP.scala 595:34]
  wire  _GEN_2807 = _GEN_145 | _GEN_2775; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2808 = _GEN_146 | _GEN_2776; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2809 = _GEN_147 | _GEN_2777; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2810 = _GEN_148 | _GEN_2778; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_2811 = 2'h0 == opidx ? 5'h5 : _GEN_2779; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2812 = 2'h1 == opidx ? 5'h5 : _GEN_2780; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2813 = 2'h2 == opidx ? 5'h5 : _GEN_2781; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2814 = 2'h3 == opidx ? 5'h5 : _GEN_2782; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_2815 = _T_122 ? _cnt_T : _GEN_2783; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_2816 = _T_122 ? _GEN_1349 : _GEN_2437; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_2817 = cnt[0] ? _GEN_2807 : _GEN_2775; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2818 = cnt[0] ? _GEN_2808 : _GEN_2776; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2819 = cnt[0] ? _GEN_2809 : _GEN_2777; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2820 = cnt[0] ? _GEN_2810 : _GEN_2778; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2821 = cnt[0] ? _GEN_2811 : _GEN_2779; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2822 = cnt[0] ? _GEN_2812 : _GEN_2780; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2823 = cnt[0] ? _GEN_2813 : _GEN_2781; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2824 = cnt[0] ? _GEN_2814 : _GEN_2782; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_2825 = cnt[0] ? _GEN_2815 : _GEN_2783; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_2826 = cnt[0] ? _GEN_2816 : _GEN_2437; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2827 = _GEN_145 | _GEN_2817; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2828 = _GEN_146 | _GEN_2818; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2829 = _GEN_147 | _GEN_2819; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_2830 = _GEN_148 | _GEN_2820; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_2831 = 2'h0 == opidx ? 5'h6 : _GEN_2821; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2832 = 2'h1 == opidx ? 5'h6 : _GEN_2822; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2833 = 2'h2 == opidx ? 5'h6 : _GEN_2823; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_2834 = 2'h3 == opidx ? 5'h6 : _GEN_2824; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_2835 = _T_122 ? _cnt_T : _GEN_2825; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_2836 = _T_122 ? _GEN_1349 : _GEN_2785; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_2837 = cnt[1] ? _GEN_2827 : _GEN_2817; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2838 = cnt[1] ? _GEN_2828 : _GEN_2818; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2839 = cnt[1] ? _GEN_2829 : _GEN_2819; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2840 = cnt[1] ? _GEN_2830 : _GEN_2820; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2841 = cnt[1] ? _GEN_2831 : _GEN_2821; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2842 = cnt[1] ? _GEN_2832 : _GEN_2822; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2843 = cnt[1] ? _GEN_2833 : _GEN_2823; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_2844 = cnt[1] ? _GEN_2834 : _GEN_2824; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_2845 = cnt[1] ? _GEN_2835 : _GEN_2825; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_2846 = cnt[1] ? _GEN_2836 : _GEN_2785; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_2847 = _GEN_145 | _GEN_2465; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_2848 = _GEN_146 | _GEN_2466; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_2849 = _GEN_147 | _GEN_2467; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_2850 = _GEN_148 | _GEN_2468; // @[NulCtrlMP.scala 377:{27,27}]
  wire [4:0] _GEN_2851 = 2'h0 == opidx ? 5'h6 : _GEN_2841; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_2852 = 2'h1 == opidx ? 5'h6 : _GEN_2842; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_2853 = 2'h2 == opidx ? 5'h6 : _GEN_2843; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_2854 = 2'h3 == opidx ? 5'h6 : _GEN_2844; // @[NulCtrlMP.scala 378:{28,28}]
  wire [63:0] _io_cpu_regacc_wdata_T_2 = {16'h0,oparg_7,oparg_6,oparg_5,oparg_4,oparg_3,oparg_2}; // @[NulCtrlMP.scala 388:53]
  wire [63:0] _GEN_2855 = 2'h0 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_2469; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_2856 = 2'h1 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_2470; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_2857 = 2'h2 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_2471; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_2858 = 2'h3 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_2472; // @[NulCtrlMP.scala 388:{30,30}]
  wire [128:0] _GEN_2859 = _T_122 ? _cnt_T : _GEN_2845; // @[NulCtrlMP.scala 389:36 390:17]
  wire  _GEN_2860 = cnt[2] ? _GEN_2847 : _GEN_2465; // @[NulCtrlMP.scala 655:22]
  wire  _GEN_2861 = cnt[2] ? _GEN_2848 : _GEN_2466; // @[NulCtrlMP.scala 655:22]
  wire  _GEN_2862 = cnt[2] ? _GEN_2849 : _GEN_2467; // @[NulCtrlMP.scala 655:22]
  wire  _GEN_2863 = cnt[2] ? _GEN_2850 : _GEN_2468; // @[NulCtrlMP.scala 655:22]
  wire [4:0] _GEN_2864 = cnt[2] ? _GEN_2851 : _GEN_2841; // @[NulCtrlMP.scala 655:22]
  wire [4:0] _GEN_2865 = cnt[2] ? _GEN_2852 : _GEN_2842; // @[NulCtrlMP.scala 655:22]
  wire [4:0] _GEN_2866 = cnt[2] ? _GEN_2853 : _GEN_2843; // @[NulCtrlMP.scala 655:22]
  wire [4:0] _GEN_2867 = cnt[2] ? _GEN_2854 : _GEN_2844; // @[NulCtrlMP.scala 655:22]
  wire [63:0] _GEN_2868 = cnt[2] ? _GEN_2855 : _GEN_2469; // @[NulCtrlMP.scala 655:22]
  wire [63:0] _GEN_2869 = cnt[2] ? _GEN_2856 : _GEN_2470; // @[NulCtrlMP.scala 655:22]
  wire [63:0] _GEN_2870 = cnt[2] ? _GEN_2857 : _GEN_2471; // @[NulCtrlMP.scala 655:22]
  wire [63:0] _GEN_2871 = cnt[2] ? _GEN_2858 : _GEN_2472; // @[NulCtrlMP.scala 655:22]
  wire [128:0] _GEN_2872 = cnt[2] ? _GEN_2859 : _GEN_2845; // @[NulCtrlMP.scala 655:22]
  wire  _GEN_2873 = _GEN_145 | _GEN_2787; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2874 = _GEN_146 | _GEN_2788; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2875 = _GEN_147 | _GEN_2789; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2876 = _GEN_148 | _GEN_2790; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2877 = 2'h0 == opidx ? 32'h34131073 : _GEN_2791; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2878 = 2'h1 == opidx ? 32'h34131073 : _GEN_2792; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2879 = 2'h2 == opidx ? 32'h34131073 : _GEN_2793; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2880 = 2'h3 == opidx ? 32'h34131073 : _GEN_2794; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2881 = _GEN_1180 ? _cnt_T : _GEN_2872; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2882 = cnt[3] ? _GEN_2873 : _GEN_2787; // @[NulCtrlMP.scala 656:22]
  wire  _GEN_2883 = cnt[3] ? _GEN_2874 : _GEN_2788; // @[NulCtrlMP.scala 656:22]
  wire  _GEN_2884 = cnt[3] ? _GEN_2875 : _GEN_2789; // @[NulCtrlMP.scala 656:22]
  wire  _GEN_2885 = cnt[3] ? _GEN_2876 : _GEN_2790; // @[NulCtrlMP.scala 656:22]
  wire [31:0] _GEN_2886 = cnt[3] ? _GEN_2877 : _GEN_2791; // @[NulCtrlMP.scala 656:22]
  wire [31:0] _GEN_2887 = cnt[3] ? _GEN_2878 : _GEN_2792; // @[NulCtrlMP.scala 656:22]
  wire [31:0] _GEN_2888 = cnt[3] ? _GEN_2879 : _GEN_2793; // @[NulCtrlMP.scala 656:22]
  wire [31:0] _GEN_2889 = cnt[3] ? _GEN_2880 : _GEN_2794; // @[NulCtrlMP.scala 656:22]
  wire [128:0] _GEN_2890 = cnt[3] ? _GEN_2881 : _GEN_2872; // @[NulCtrlMP.scala 656:22]
  wire  _GEN_2891 = _GEN_145 | _GEN_2882; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2892 = _GEN_146 | _GEN_2883; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2893 = _GEN_147 | _GEN_2884; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2894 = _GEN_148 | _GEN_2885; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2895 = 2'h0 == opidx ? 32'h300293 : _GEN_2886; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2896 = 2'h1 == opidx ? 32'h300293 : _GEN_2887; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2897 = 2'h2 == opidx ? 32'h300293 : _GEN_2888; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2898 = 2'h3 == opidx ? 32'h300293 : _GEN_2889; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2899 = _GEN_1180 ? _cnt_T : _GEN_2890; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2900 = cnt[4] ? _GEN_2891 : _GEN_2882; // @[NulCtrlMP.scala 658:22]
  wire  _GEN_2901 = cnt[4] ? _GEN_2892 : _GEN_2883; // @[NulCtrlMP.scala 658:22]
  wire  _GEN_2902 = cnt[4] ? _GEN_2893 : _GEN_2884; // @[NulCtrlMP.scala 658:22]
  wire  _GEN_2903 = cnt[4] ? _GEN_2894 : _GEN_2885; // @[NulCtrlMP.scala 658:22]
  wire [31:0] _GEN_2904 = cnt[4] ? _GEN_2895 : _GEN_2886; // @[NulCtrlMP.scala 658:22]
  wire [31:0] _GEN_2905 = cnt[4] ? _GEN_2896 : _GEN_2887; // @[NulCtrlMP.scala 658:22]
  wire [31:0] _GEN_2906 = cnt[4] ? _GEN_2897 : _GEN_2888; // @[NulCtrlMP.scala 658:22]
  wire [31:0] _GEN_2907 = cnt[4] ? _GEN_2898 : _GEN_2889; // @[NulCtrlMP.scala 658:22]
  wire [128:0] _GEN_2908 = cnt[4] ? _GEN_2899 : _GEN_2890; // @[NulCtrlMP.scala 658:22]
  wire  _GEN_2909 = _GEN_145 | _GEN_2900; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2910 = _GEN_146 | _GEN_2901; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2911 = _GEN_147 | _GEN_2902; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2912 = _GEN_148 | _GEN_2903; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2913 = 2'h0 == opidx ? 32'hb29293 : _GEN_2904; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2914 = 2'h1 == opidx ? 32'hb29293 : _GEN_2905; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2915 = 2'h2 == opidx ? 32'hb29293 : _GEN_2906; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2916 = 2'h3 == opidx ? 32'hb29293 : _GEN_2907; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2917 = _GEN_1180 ? _cnt_T : _GEN_2908; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2918 = cnt[5] ? _GEN_2909 : _GEN_2900; // @[NulCtrlMP.scala 659:22]
  wire  _GEN_2919 = cnt[5] ? _GEN_2910 : _GEN_2901; // @[NulCtrlMP.scala 659:22]
  wire  _GEN_2920 = cnt[5] ? _GEN_2911 : _GEN_2902; // @[NulCtrlMP.scala 659:22]
  wire  _GEN_2921 = cnt[5] ? _GEN_2912 : _GEN_2903; // @[NulCtrlMP.scala 659:22]
  wire [31:0] _GEN_2922 = cnt[5] ? _GEN_2913 : _GEN_2904; // @[NulCtrlMP.scala 659:22]
  wire [31:0] _GEN_2923 = cnt[5] ? _GEN_2914 : _GEN_2905; // @[NulCtrlMP.scala 659:22]
  wire [31:0] _GEN_2924 = cnt[5] ? _GEN_2915 : _GEN_2906; // @[NulCtrlMP.scala 659:22]
  wire [31:0] _GEN_2925 = cnt[5] ? _GEN_2916 : _GEN_2907; // @[NulCtrlMP.scala 659:22]
  wire [128:0] _GEN_2926 = cnt[5] ? _GEN_2917 : _GEN_2908; // @[NulCtrlMP.scala 659:22]
  wire  _GEN_2927 = _GEN_145 | _GEN_2918; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2928 = _GEN_146 | _GEN_2919; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2929 = _GEN_147 | _GEN_2920; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2930 = _GEN_148 | _GEN_2921; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2931 = 2'h0 == opidx ? 32'h3002b073 : _GEN_2922; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2932 = 2'h1 == opidx ? 32'h3002b073 : _GEN_2923; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2933 = 2'h2 == opidx ? 32'h3002b073 : _GEN_2924; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2934 = 2'h3 == opidx ? 32'h3002b073 : _GEN_2925; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2935 = _GEN_1180 ? _cnt_T : _GEN_2926; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2936 = cnt[6] ? _GEN_2927 : _GEN_2918; // @[NulCtrlMP.scala 660:22]
  wire  _GEN_2937 = cnt[6] ? _GEN_2928 : _GEN_2919; // @[NulCtrlMP.scala 660:22]
  wire  _GEN_2938 = cnt[6] ? _GEN_2929 : _GEN_2920; // @[NulCtrlMP.scala 660:22]
  wire  _GEN_2939 = cnt[6] ? _GEN_2930 : _GEN_2921; // @[NulCtrlMP.scala 660:22]
  wire [31:0] _GEN_2940 = cnt[6] ? _GEN_2931 : _GEN_2922; // @[NulCtrlMP.scala 660:22]
  wire [31:0] _GEN_2941 = cnt[6] ? _GEN_2932 : _GEN_2923; // @[NulCtrlMP.scala 660:22]
  wire [31:0] _GEN_2942 = cnt[6] ? _GEN_2933 : _GEN_2924; // @[NulCtrlMP.scala 660:22]
  wire [31:0] _GEN_2943 = cnt[6] ? _GEN_2934 : _GEN_2925; // @[NulCtrlMP.scala 660:22]
  wire [128:0] _GEN_2944 = cnt[6] ? _GEN_2935 : _GEN_2926; // @[NulCtrlMP.scala 660:22]
  wire  _GEN_2945 = _GEN_145 | _GEN_2936; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2946 = _GEN_146 | _GEN_2937; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2947 = _GEN_147 | _GEN_2938; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2948 = _GEN_148 | _GEN_2939; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2949 = 2'h0 == opidx ? 32'h22b7 : _GEN_2940; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2950 = 2'h1 == opidx ? 32'h22b7 : _GEN_2941; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2951 = 2'h2 == opidx ? 32'h22b7 : _GEN_2942; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2952 = 2'h3 == opidx ? 32'h22b7 : _GEN_2943; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2953 = _GEN_1180 ? _cnt_T : _GEN_2944; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2954 = cnt[7] ? _GEN_2945 : _GEN_2936; // @[NulCtrlMP.scala 661:22]
  wire  _GEN_2955 = cnt[7] ? _GEN_2946 : _GEN_2937; // @[NulCtrlMP.scala 661:22]
  wire  _GEN_2956 = cnt[7] ? _GEN_2947 : _GEN_2938; // @[NulCtrlMP.scala 661:22]
  wire  _GEN_2957 = cnt[7] ? _GEN_2948 : _GEN_2939; // @[NulCtrlMP.scala 661:22]
  wire [31:0] _GEN_2958 = cnt[7] ? _GEN_2949 : _GEN_2940; // @[NulCtrlMP.scala 661:22]
  wire [31:0] _GEN_2959 = cnt[7] ? _GEN_2950 : _GEN_2941; // @[NulCtrlMP.scala 661:22]
  wire [31:0] _GEN_2960 = cnt[7] ? _GEN_2951 : _GEN_2942; // @[NulCtrlMP.scala 661:22]
  wire [31:0] _GEN_2961 = cnt[7] ? _GEN_2952 : _GEN_2943; // @[NulCtrlMP.scala 661:22]
  wire [128:0] _GEN_2962 = cnt[7] ? _GEN_2953 : _GEN_2944; // @[NulCtrlMP.scala 661:22]
  wire  _GEN_2963 = _GEN_145 | _GEN_2954; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2964 = _GEN_146 | _GEN_2955; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2965 = _GEN_147 | _GEN_2956; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2966 = _GEN_148 | _GEN_2957; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2967 = 2'h0 == opidx ? 32'h3002a073 : _GEN_2958; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2968 = 2'h1 == opidx ? 32'h3002a073 : _GEN_2959; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2969 = 2'h2 == opidx ? 32'h3002a073 : _GEN_2960; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2970 = 2'h3 == opidx ? 32'h3002a073 : _GEN_2961; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2971 = _GEN_1180 ? _cnt_T : _GEN_2962; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2972 = cnt[8] ? _GEN_2963 : _GEN_2954; // @[NulCtrlMP.scala 668:22]
  wire  _GEN_2973 = cnt[8] ? _GEN_2964 : _GEN_2955; // @[NulCtrlMP.scala 668:22]
  wire  _GEN_2974 = cnt[8] ? _GEN_2965 : _GEN_2956; // @[NulCtrlMP.scala 668:22]
  wire  _GEN_2975 = cnt[8] ? _GEN_2966 : _GEN_2957; // @[NulCtrlMP.scala 668:22]
  wire [31:0] _GEN_2976 = cnt[8] ? _GEN_2967 : _GEN_2958; // @[NulCtrlMP.scala 668:22]
  wire [31:0] _GEN_2977 = cnt[8] ? _GEN_2968 : _GEN_2959; // @[NulCtrlMP.scala 668:22]
  wire [31:0] _GEN_2978 = cnt[8] ? _GEN_2969 : _GEN_2960; // @[NulCtrlMP.scala 668:22]
  wire [31:0] _GEN_2979 = cnt[8] ? _GEN_2970 : _GEN_2961; // @[NulCtrlMP.scala 668:22]
  wire [128:0] _GEN_2980 = cnt[8] ? _GEN_2971 : _GEN_2962; // @[NulCtrlMP.scala 668:22]
  wire  _GEN_2981 = _GEN_145 | _GEN_2972; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2982 = _GEN_146 | _GEN_2973; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2983 = _GEN_147 | _GEN_2974; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_2984 = _GEN_148 | _GEN_2975; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_2985 = 2'h0 == opidx ? 32'h301073 : _GEN_2976; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2986 = 2'h1 == opidx ? 32'h301073 : _GEN_2977; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2987 = 2'h2 == opidx ? 32'h301073 : _GEN_2978; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_2988 = 2'h3 == opidx ? 32'h301073 : _GEN_2979; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_2989 = _GEN_1180 ? _cnt_T : _GEN_2980; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_2990 = cnt[9] ? _GEN_2981 : _GEN_2972; // @[NulCtrlMP.scala 675:22]
  wire  _GEN_2991 = cnt[9] ? _GEN_2982 : _GEN_2973; // @[NulCtrlMP.scala 675:22]
  wire  _GEN_2992 = cnt[9] ? _GEN_2983 : _GEN_2974; // @[NulCtrlMP.scala 675:22]
  wire  _GEN_2993 = cnt[9] ? _GEN_2984 : _GEN_2975; // @[NulCtrlMP.scala 675:22]
  wire [31:0] _GEN_2994 = cnt[9] ? _GEN_2985 : _GEN_2976; // @[NulCtrlMP.scala 675:22]
  wire [31:0] _GEN_2995 = cnt[9] ? _GEN_2986 : _GEN_2977; // @[NulCtrlMP.scala 675:22]
  wire [31:0] _GEN_2996 = cnt[9] ? _GEN_2987 : _GEN_2978; // @[NulCtrlMP.scala 675:22]
  wire [31:0] _GEN_2997 = cnt[9] ? _GEN_2988 : _GEN_2979; // @[NulCtrlMP.scala 675:22]
  wire [128:0] _GEN_2998 = cnt[9] ? _GEN_2989 : _GEN_2980; // @[NulCtrlMP.scala 675:22]
  wire  _GEN_2999 = _GEN_145 | _GEN_2990; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3000 = _GEN_146 | _GEN_2991; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3001 = _GEN_147 | _GEN_2992; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3002 = _GEN_148 | _GEN_2993; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3003 = 2'h0 == opidx ? 32'h330000f : _GEN_2994; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3004 = 2'h1 == opidx ? 32'h330000f : _GEN_2995; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3005 = 2'h2 == opidx ? 32'h330000f : _GEN_2996; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3006 = 2'h3 == opidx ? 32'h330000f : _GEN_2997; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3007 = _GEN_1180 ? _cnt_T : _GEN_2998; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3008 = cnt[10] ? _GEN_2999 : _GEN_2990; // @[NulCtrlMP.scala 682:23]
  wire  _GEN_3009 = cnt[10] ? _GEN_3000 : _GEN_2991; // @[NulCtrlMP.scala 682:23]
  wire  _GEN_3010 = cnt[10] ? _GEN_3001 : _GEN_2992; // @[NulCtrlMP.scala 682:23]
  wire  _GEN_3011 = cnt[10] ? _GEN_3002 : _GEN_2993; // @[NulCtrlMP.scala 682:23]
  wire [31:0] _GEN_3012 = cnt[10] ? _GEN_3003 : _GEN_2994; // @[NulCtrlMP.scala 682:23]
  wire [31:0] _GEN_3013 = cnt[10] ? _GEN_3004 : _GEN_2995; // @[NulCtrlMP.scala 682:23]
  wire [31:0] _GEN_3014 = cnt[10] ? _GEN_3005 : _GEN_2996; // @[NulCtrlMP.scala 682:23]
  wire [31:0] _GEN_3015 = cnt[10] ? _GEN_3006 : _GEN_2997; // @[NulCtrlMP.scala 682:23]
  wire [128:0] _GEN_3016 = cnt[10] ? _GEN_3007 : _GEN_2998; // @[NulCtrlMP.scala 682:23]
  wire  _GEN_3017 = _GEN_145 | _GEN_2795; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3018 = _GEN_146 | _GEN_2796; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3019 = _GEN_147 | _GEN_2797; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3020 = _GEN_148 | _GEN_2798; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_3021 = ~_GEN_1252 ? _cnt_T : _GEN_3016; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_3022 = cnt[11] ? _GEN_3017 : _GEN_2795; // @[NulCtrlMP.scala 683:23]
  wire  _GEN_3023 = cnt[11] ? _GEN_3018 : _GEN_2796; // @[NulCtrlMP.scala 683:23]
  wire  _GEN_3024 = cnt[11] ? _GEN_3019 : _GEN_2797; // @[NulCtrlMP.scala 683:23]
  wire  _GEN_3025 = cnt[11] ? _GEN_3020 : _GEN_2798; // @[NulCtrlMP.scala 683:23]
  wire [128:0] _GEN_3026 = cnt[11] ? _GEN_3021 : _GEN_3016; // @[NulCtrlMP.scala 683:23]
  wire  _GEN_3027 = _GEN_145 | _GEN_2860; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3028 = _GEN_146 | _GEN_2861; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3029 = _GEN_147 | _GEN_2862; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3030 = _GEN_148 | _GEN_2863; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_3031 = 2'h0 == opidx ? 5'h5 : _GEN_2864; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3032 = 2'h1 == opidx ? 5'h5 : _GEN_2865; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3033 = 2'h2 == opidx ? 5'h5 : _GEN_2866; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3034 = 2'h3 == opidx ? 5'h5 : _GEN_2867; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_3035 = 2'h0 == opidx ? regback_0 : _GEN_2868; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3036 = 2'h1 == opidx ? regback_0 : _GEN_2869; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3037 = 2'h2 == opidx ? regback_0 : _GEN_2870; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3038 = 2'h3 == opidx ? regback_0 : _GEN_2871; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_3039 = ~_GEN_1128 ? _cnt_T : _GEN_3026; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_3040 = cnt[12] ? _GEN_3027 : _GEN_2860; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3041 = cnt[12] ? _GEN_3028 : _GEN_2861; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3042 = cnt[12] ? _GEN_3029 : _GEN_2862; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3043 = cnt[12] ? _GEN_3030 : _GEN_2863; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3044 = cnt[12] ? _GEN_3031 : _GEN_2864; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3045 = cnt[12] ? _GEN_3032 : _GEN_2865; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3046 = cnt[12] ? _GEN_3033 : _GEN_2866; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3047 = cnt[12] ? _GEN_3034 : _GEN_2867; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3048 = cnt[12] ? _GEN_3035 : _GEN_2868; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3049 = cnt[12] ? _GEN_3036 : _GEN_2869; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3050 = cnt[12] ? _GEN_3037 : _GEN_2870; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3051 = cnt[12] ? _GEN_3038 : _GEN_2871; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3052 = cnt[12] ? _GEN_3039 : _GEN_3026; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3053 = _GEN_145 | _GEN_3040; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3054 = _GEN_146 | _GEN_3041; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3055 = _GEN_147 | _GEN_3042; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3056 = _GEN_148 | _GEN_3043; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_3057 = 2'h0 == opidx ? 5'h6 : _GEN_3044; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3058 = 2'h1 == opidx ? 5'h6 : _GEN_3045; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3059 = 2'h2 == opidx ? 5'h6 : _GEN_3046; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3060 = 2'h3 == opidx ? 5'h6 : _GEN_3047; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_3061 = 2'h0 == opidx ? regback_1 : _GEN_3048; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3062 = 2'h1 == opidx ? regback_1 : _GEN_3049; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3063 = 2'h2 == opidx ? regback_1 : _GEN_3050; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3064 = 2'h3 == opidx ? regback_1 : _GEN_3051; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_3065 = ~_GEN_1128 ? _cnt_T : _GEN_3052; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_3066 = cnt[13] ? _GEN_3053 : _GEN_3040; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3067 = cnt[13] ? _GEN_3054 : _GEN_3041; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3068 = cnt[13] ? _GEN_3055 : _GEN_3042; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3069 = cnt[13] ? _GEN_3056 : _GEN_3043; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3070 = cnt[13] ? _GEN_3057 : _GEN_3044; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3071 = cnt[13] ? _GEN_3058 : _GEN_3045; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3072 = cnt[13] ? _GEN_3059 : _GEN_3046; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3073 = cnt[13] ? _GEN_3060 : _GEN_3047; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3074 = cnt[13] ? _GEN_3061 : _GEN_3048; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3075 = cnt[13] ? _GEN_3062 : _GEN_3049; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3076 = cnt[13] ? _GEN_3063 : _GEN_3050; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3077 = cnt[13] ? _GEN_3064 : _GEN_3051; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3078 = cnt[13] ? _GEN_3065 : _GEN_3052; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3079 = _GEN_145 | _GEN_2799; // @[NulCtrlMP.scala 686:{35,35}]
  wire  _GEN_3080 = _GEN_146 | _GEN_2800; // @[NulCtrlMP.scala 686:{35,35}]
  wire  _GEN_3081 = _GEN_147 | _GEN_2801; // @[NulCtrlMP.scala 686:{35,35}]
  wire  _GEN_3082 = _GEN_148 | _GEN_2802; // @[NulCtrlMP.scala 686:{35,35}]
  wire  _GEN_3083 = _GEN_145 | _GEN_3008; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3084 = _GEN_146 | _GEN_3009; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3085 = _GEN_147 | _GEN_3010; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3086 = _GEN_148 | _GEN_3011; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3087 = 2'h0 == opidx ? 32'h30200073 : _GEN_3012; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3088 = 2'h1 == opidx ? 32'h30200073 : _GEN_3013; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3089 = 2'h2 == opidx ? 32'h30200073 : _GEN_3014; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3090 = 2'h3 == opidx ? 32'h30200073 : _GEN_3015; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3091 = _GEN_1180 ? _cnt_T : _GEN_3078; // @[NulCtrlMP.scala 396:36 397:17]
  wire [1:0] _GEN_3092 = 2'h0 == opidx ? 2'h3 : _GEN_2803; // @[NulCtrlMP.scala 689:{34,34}]
  wire [1:0] _GEN_3093 = 2'h1 == opidx ? 2'h3 : _GEN_2804; // @[NulCtrlMP.scala 689:{34,34}]
  wire [1:0] _GEN_3094 = 2'h2 == opidx ? 2'h3 : _GEN_2805; // @[NulCtrlMP.scala 689:{34,34}]
  wire [1:0] _GEN_3095 = 2'h3 == opidx ? 2'h3 : _GEN_2806; // @[NulCtrlMP.scala 689:{34,34}]
  wire  _GEN_3100 = cnt[14] ? _GEN_3079 : _GEN_2799; // @[NulCtrlMP.scala 685:23]
  wire  _GEN_3101 = cnt[14] ? _GEN_3080 : _GEN_2800; // @[NulCtrlMP.scala 685:23]
  wire  _GEN_3102 = cnt[14] ? _GEN_3081 : _GEN_2801; // @[NulCtrlMP.scala 685:23]
  wire  _GEN_3103 = cnt[14] ? _GEN_3082 : _GEN_2802; // @[NulCtrlMP.scala 685:23]
  wire  _GEN_3104 = cnt[14] ? _GEN_3083 : _GEN_3008; // @[NulCtrlMP.scala 685:23]
  wire  _GEN_3105 = cnt[14] ? _GEN_3084 : _GEN_3009; // @[NulCtrlMP.scala 685:23]
  wire  _GEN_3106 = cnt[14] ? _GEN_3085 : _GEN_3010; // @[NulCtrlMP.scala 685:23]
  wire  _GEN_3107 = cnt[14] ? _GEN_3086 : _GEN_3011; // @[NulCtrlMP.scala 685:23]
  wire [31:0] _GEN_3108 = cnt[14] ? _GEN_3087 : _GEN_3012; // @[NulCtrlMP.scala 685:23]
  wire [31:0] _GEN_3109 = cnt[14] ? _GEN_3088 : _GEN_3013; // @[NulCtrlMP.scala 685:23]
  wire [31:0] _GEN_3110 = cnt[14] ? _GEN_3089 : _GEN_3014; // @[NulCtrlMP.scala 685:23]
  wire [31:0] _GEN_3111 = cnt[14] ? _GEN_3090 : _GEN_3015; // @[NulCtrlMP.scala 685:23]
  wire [128:0] _GEN_3112 = cnt[14] ? _GEN_3091 : _GEN_3078; // @[NulCtrlMP.scala 685:23]
  wire  _GEN_3117 = _GEN_145 | _GEN_3022; // @[NulCtrlMP.scala 693:{34,34}]
  wire  _GEN_3118 = _GEN_146 | _GEN_3023; // @[NulCtrlMP.scala 693:{34,34}]
  wire  _GEN_3119 = _GEN_147 | _GEN_3024; // @[NulCtrlMP.scala 693:{34,34}]
  wire  _GEN_3120 = _GEN_148 | _GEN_3025; // @[NulCtrlMP.scala 693:{34,34}]
  wire  _GEN_3121 = cnt[15] ? _GEN_3117 : _GEN_3022; // @[NulCtrlMP.scala 692:23]
  wire  _GEN_3122 = cnt[15] ? _GEN_3118 : _GEN_3023; // @[NulCtrlMP.scala 692:23]
  wire  _GEN_3123 = cnt[15] ? _GEN_3119 : _GEN_3024; // @[NulCtrlMP.scala 692:23]
  wire  _GEN_3124 = cnt[15] ? _GEN_3120 : _GEN_3025; // @[NulCtrlMP.scala 692:23]
  wire [128:0] _GEN_3125 = cnt[15] ? _cnt_T : _GEN_3112; // @[NulCtrlMP.scala 692:23 694:17]
  wire [128:0] _GEN_3126 = cnt[16] ? 129'h1 : _GEN_3125; // @[NulCtrlMP.scala 696:23 697:17]
  wire [4:0] _GEN_3127 = cnt[16] ? 5'h5 : _GEN_2786; // @[NulCtrlMP.scala 696:23 698:19]
  wire  _GEN_3128 = state == 5'hb ? _GEN_2837 : _GEN_2775; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3129 = state == 5'hb ? _GEN_2838 : _GEN_2776; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3130 = state == 5'hb ? _GEN_2839 : _GEN_2777; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3131 = state == 5'hb ? _GEN_2840 : _GEN_2778; // @[NulCtrlMP.scala 653:33]
  wire [4:0] _GEN_3132 = state == 5'hb ? _GEN_3070 : _GEN_2779; // @[NulCtrlMP.scala 653:33]
  wire [4:0] _GEN_3133 = state == 5'hb ? _GEN_3071 : _GEN_2780; // @[NulCtrlMP.scala 653:33]
  wire [4:0] _GEN_3134 = state == 5'hb ? _GEN_3072 : _GEN_2781; // @[NulCtrlMP.scala 653:33]
  wire [4:0] _GEN_3135 = state == 5'hb ? _GEN_3073 : _GEN_2782; // @[NulCtrlMP.scala 653:33]
  wire [128:0] _GEN_3136 = state == 5'hb ? _GEN_3126 : _GEN_2783; // @[NulCtrlMP.scala 653:33]
  wire [63:0] _GEN_3137 = state == 5'hb ? _GEN_2826 : _GEN_2437; // @[NulCtrlMP.scala 653:33]
  wire [63:0] _GEN_3138 = state == 5'hb ? _GEN_2846 : _GEN_2785; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3139 = state == 5'hb ? _GEN_3066 : _GEN_2465; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3140 = state == 5'hb ? _GEN_3067 : _GEN_2466; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3141 = state == 5'hb ? _GEN_3068 : _GEN_2467; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3142 = state == 5'hb ? _GEN_3069 : _GEN_2468; // @[NulCtrlMP.scala 653:33]
  wire [63:0] _GEN_3143 = state == 5'hb ? _GEN_3074 : _GEN_2469; // @[NulCtrlMP.scala 653:33]
  wire [63:0] _GEN_3144 = state == 5'hb ? _GEN_3075 : _GEN_2470; // @[NulCtrlMP.scala 653:33]
  wire [63:0] _GEN_3145 = state == 5'hb ? _GEN_3076 : _GEN_2471; // @[NulCtrlMP.scala 653:33]
  wire [63:0] _GEN_3146 = state == 5'hb ? _GEN_3077 : _GEN_2472; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3147 = state == 5'hb ? _GEN_3104 : _GEN_2787; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3148 = state == 5'hb ? _GEN_3105 : _GEN_2788; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3149 = state == 5'hb ? _GEN_3106 : _GEN_2789; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3150 = state == 5'hb ? _GEN_3107 : _GEN_2790; // @[NulCtrlMP.scala 653:33]
  wire [31:0] _GEN_3151 = state == 5'hb ? _GEN_3108 : _GEN_2791; // @[NulCtrlMP.scala 653:33]
  wire [31:0] _GEN_3152 = state == 5'hb ? _GEN_3109 : _GEN_2792; // @[NulCtrlMP.scala 653:33]
  wire [31:0] _GEN_3153 = state == 5'hb ? _GEN_3110 : _GEN_2793; // @[NulCtrlMP.scala 653:33]
  wire [31:0] _GEN_3154 = state == 5'hb ? _GEN_3111 : _GEN_2794; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3155 = state == 5'hb ? _GEN_3121 : _GEN_2795; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3156 = state == 5'hb ? _GEN_3122 : _GEN_2796; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3157 = state == 5'hb ? _GEN_3123 : _GEN_2797; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3158 = state == 5'hb ? _GEN_3124 : _GEN_2798; // @[NulCtrlMP.scala 653:33]
  wire [4:0] _GEN_3167 = state == 5'hb ? _GEN_3127 : _GEN_2786; // @[NulCtrlMP.scala 653:33]
  wire  _GEN_3168 = _GEN_145 | _GEN_3128; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3169 = _GEN_146 | _GEN_3129; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3170 = _GEN_147 | _GEN_3130; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3171 = _GEN_148 | _GEN_3131; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_3172 = 2'h0 == opidx ? 5'h5 : _GEN_3132; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3173 = 2'h1 == opidx ? 5'h5 : _GEN_3133; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3174 = 2'h2 == opidx ? 5'h5 : _GEN_3134; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3175 = 2'h3 == opidx ? 5'h5 : _GEN_3135; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_3176 = _T_122 ? _cnt_T : _GEN_3136; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_3177 = _T_122 ? _GEN_1349 : _GEN_3137; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_3178 = cnt[0] ? _GEN_3168 : _GEN_3128; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3179 = cnt[0] ? _GEN_3169 : _GEN_3129; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3180 = cnt[0] ? _GEN_3170 : _GEN_3130; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3181 = cnt[0] ? _GEN_3171 : _GEN_3131; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3182 = cnt[0] ? _GEN_3172 : _GEN_3132; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3183 = cnt[0] ? _GEN_3173 : _GEN_3133; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3184 = cnt[0] ? _GEN_3174 : _GEN_3134; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3185 = cnt[0] ? _GEN_3175 : _GEN_3135; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_3186 = cnt[0] ? _GEN_3176 : _GEN_3136; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_3187 = cnt[0] ? _GEN_3177 : _GEN_3137; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3188 = _GEN_145 | _GEN_3178; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3189 = _GEN_146 | _GEN_3179; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3190 = _GEN_147 | _GEN_3180; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3191 = _GEN_148 | _GEN_3181; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_3192 = 2'h0 == opidx ? 5'h6 : _GEN_3182; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3193 = 2'h1 == opidx ? 5'h6 : _GEN_3183; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3194 = 2'h2 == opidx ? 5'h6 : _GEN_3184; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3195 = 2'h3 == opidx ? 5'h6 : _GEN_3185; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_3196 = _T_122 ? _cnt_T : _GEN_3186; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_3197 = _T_122 ? _GEN_1349 : _GEN_3138; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_3198 = cnt[1] ? _GEN_3188 : _GEN_3178; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3199 = cnt[1] ? _GEN_3189 : _GEN_3179; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3200 = cnt[1] ? _GEN_3190 : _GEN_3180; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3201 = cnt[1] ? _GEN_3191 : _GEN_3181; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3202 = cnt[1] ? _GEN_3192 : _GEN_3182; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3203 = cnt[1] ? _GEN_3193 : _GEN_3183; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3204 = cnt[1] ? _GEN_3194 : _GEN_3184; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3205 = cnt[1] ? _GEN_3195 : _GEN_3185; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_3206 = cnt[1] ? _GEN_3196 : _GEN_3186; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_3207 = cnt[1] ? _GEN_3197 : _GEN_3138; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3208 = _GEN_145 | _GEN_3139; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3209 = _GEN_146 | _GEN_3140; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3210 = _GEN_147 | _GEN_3141; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3211 = _GEN_148 | _GEN_3142; // @[NulCtrlMP.scala 377:{27,27}]
  wire [4:0] _GEN_3212 = 2'h0 == opidx ? 5'h5 : _GEN_3202; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3213 = 2'h1 == opidx ? 5'h5 : _GEN_3203; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3214 = 2'h2 == opidx ? 5'h5 : _GEN_3204; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3215 = 2'h3 == opidx ? 5'h5 : _GEN_3205; // @[NulCtrlMP.scala 378:{28,28}]
  wire [63:0] _GEN_3216 = 2'h0 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_3143; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3217 = 2'h1 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_3144; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3218 = 2'h2 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_3145; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3219 = 2'h3 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_3146; // @[NulCtrlMP.scala 388:{30,30}]
  wire [128:0] _GEN_3220 = _T_122 ? _cnt_T : _GEN_3206; // @[NulCtrlMP.scala 389:36 390:17]
  wire  _GEN_3221 = cnt[2] ? _GEN_3208 : _GEN_3139; // @[NulCtrlMP.scala 704:22]
  wire  _GEN_3222 = cnt[2] ? _GEN_3209 : _GEN_3140; // @[NulCtrlMP.scala 704:22]
  wire  _GEN_3223 = cnt[2] ? _GEN_3210 : _GEN_3141; // @[NulCtrlMP.scala 704:22]
  wire  _GEN_3224 = cnt[2] ? _GEN_3211 : _GEN_3142; // @[NulCtrlMP.scala 704:22]
  wire [4:0] _GEN_3225 = cnt[2] ? _GEN_3212 : _GEN_3202; // @[NulCtrlMP.scala 704:22]
  wire [4:0] _GEN_3226 = cnt[2] ? _GEN_3213 : _GEN_3203; // @[NulCtrlMP.scala 704:22]
  wire [4:0] _GEN_3227 = cnt[2] ? _GEN_3214 : _GEN_3204; // @[NulCtrlMP.scala 704:22]
  wire [4:0] _GEN_3228 = cnt[2] ? _GEN_3215 : _GEN_3205; // @[NulCtrlMP.scala 704:22]
  wire [63:0] _GEN_3229 = cnt[2] ? _GEN_3216 : _GEN_3143; // @[NulCtrlMP.scala 704:22]
  wire [63:0] _GEN_3230 = cnt[2] ? _GEN_3217 : _GEN_3144; // @[NulCtrlMP.scala 704:22]
  wire [63:0] _GEN_3231 = cnt[2] ? _GEN_3218 : _GEN_3145; // @[NulCtrlMP.scala 704:22]
  wire [63:0] _GEN_3232 = cnt[2] ? _GEN_3219 : _GEN_3146; // @[NulCtrlMP.scala 704:22]
  wire [128:0] _GEN_3233 = cnt[2] ? _GEN_3220 : _GEN_3206; // @[NulCtrlMP.scala 704:22]
  wire  _GEN_3234 = _GEN_145 | _GEN_3147; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3235 = _GEN_146 | _GEN_3148; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3236 = _GEN_147 | _GEN_3149; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3237 = _GEN_148 | _GEN_3150; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3238 = 2'h0 == opidx ? 32'h2b303 : _GEN_3151; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3239 = 2'h1 == opidx ? 32'h2b303 : _GEN_3152; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3240 = 2'h2 == opidx ? 32'h2b303 : _GEN_3153; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3241 = 2'h3 == opidx ? 32'h2b303 : _GEN_3154; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3242 = _GEN_1180 ? _cnt_T : _GEN_3233; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3243 = cnt[3] ? _GEN_3234 : _GEN_3147; // @[NulCtrlMP.scala 705:22]
  wire  _GEN_3244 = cnt[3] ? _GEN_3235 : _GEN_3148; // @[NulCtrlMP.scala 705:22]
  wire  _GEN_3245 = cnt[3] ? _GEN_3236 : _GEN_3149; // @[NulCtrlMP.scala 705:22]
  wire  _GEN_3246 = cnt[3] ? _GEN_3237 : _GEN_3150; // @[NulCtrlMP.scala 705:22]
  wire [31:0] _GEN_3247 = cnt[3] ? _GEN_3238 : _GEN_3151; // @[NulCtrlMP.scala 705:22]
  wire [31:0] _GEN_3248 = cnt[3] ? _GEN_3239 : _GEN_3152; // @[NulCtrlMP.scala 705:22]
  wire [31:0] _GEN_3249 = cnt[3] ? _GEN_3240 : _GEN_3153; // @[NulCtrlMP.scala 705:22]
  wire [31:0] _GEN_3250 = cnt[3] ? _GEN_3241 : _GEN_3154; // @[NulCtrlMP.scala 705:22]
  wire [128:0] _GEN_3251 = cnt[3] ? _GEN_3242 : _GEN_3233; // @[NulCtrlMP.scala 705:22]
  wire  _GEN_3252 = _GEN_145 | _GEN_3243; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3253 = _GEN_146 | _GEN_3244; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3254 = _GEN_147 | _GEN_3245; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3255 = _GEN_148 | _GEN_3246; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3256 = 2'h0 == opidx ? 32'h330000f : _GEN_3247; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3257 = 2'h1 == opidx ? 32'h330000f : _GEN_3248; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3258 = 2'h2 == opidx ? 32'h330000f : _GEN_3249; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3259 = 2'h3 == opidx ? 32'h330000f : _GEN_3250; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3260 = _GEN_1180 ? _cnt_T : _GEN_3251; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3261 = cnt[4] ? _GEN_3252 : _GEN_3243; // @[NulCtrlMP.scala 706:22]
  wire  _GEN_3262 = cnt[4] ? _GEN_3253 : _GEN_3244; // @[NulCtrlMP.scala 706:22]
  wire  _GEN_3263 = cnt[4] ? _GEN_3254 : _GEN_3245; // @[NulCtrlMP.scala 706:22]
  wire  _GEN_3264 = cnt[4] ? _GEN_3255 : _GEN_3246; // @[NulCtrlMP.scala 706:22]
  wire [31:0] _GEN_3265 = cnt[4] ? _GEN_3256 : _GEN_3247; // @[NulCtrlMP.scala 706:22]
  wire [31:0] _GEN_3266 = cnt[4] ? _GEN_3257 : _GEN_3248; // @[NulCtrlMP.scala 706:22]
  wire [31:0] _GEN_3267 = cnt[4] ? _GEN_3258 : _GEN_3249; // @[NulCtrlMP.scala 706:22]
  wire [31:0] _GEN_3268 = cnt[4] ? _GEN_3259 : _GEN_3250; // @[NulCtrlMP.scala 706:22]
  wire [128:0] _GEN_3269 = cnt[4] ? _GEN_3260 : _GEN_3251; // @[NulCtrlMP.scala 706:22]
  wire  _GEN_3270 = _GEN_145 | _GEN_3155; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3271 = _GEN_146 | _GEN_3156; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3272 = _GEN_147 | _GEN_3157; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3273 = _GEN_148 | _GEN_3158; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_3274 = ~_GEN_1252 ? _cnt_T : _GEN_3269; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_3275 = cnt[5] ? _GEN_3270 : _GEN_3155; // @[NulCtrlMP.scala 707:22]
  wire  _GEN_3276 = cnt[5] ? _GEN_3271 : _GEN_3156; // @[NulCtrlMP.scala 707:22]
  wire  _GEN_3277 = cnt[5] ? _GEN_3272 : _GEN_3157; // @[NulCtrlMP.scala 707:22]
  wire  _GEN_3278 = cnt[5] ? _GEN_3273 : _GEN_3158; // @[NulCtrlMP.scala 707:22]
  wire [128:0] _GEN_3279 = cnt[5] ? _GEN_3274 : _GEN_3269; // @[NulCtrlMP.scala 707:22]
  wire  _GEN_3280 = _GEN_145 | _GEN_3198; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_3281 = _GEN_146 | _GEN_3199; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_3282 = _GEN_147 | _GEN_3200; // @[NulCtrlMP.scala 359:{27,27}]
  wire  _GEN_3283 = _GEN_148 | _GEN_3201; // @[NulCtrlMP.scala 359:{27,27}]
  wire [4:0] _GEN_3284 = 2'h0 == opidx ? 5'h6 : _GEN_3225; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_3285 = 2'h1 == opidx ? 5'h6 : _GEN_3226; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_3286 = 2'h2 == opidx ? 5'h6 : _GEN_3227; // @[NulCtrlMP.scala 360:{28,28}]
  wire [4:0] _GEN_3287 = 2'h3 == opidx ? 5'h6 : _GEN_3228; // @[NulCtrlMP.scala 360:{28,28}]
  wire [128:0] _GEN_3288 = _T_122 ? _cnt_T : _GEN_3279; // @[NulCtrlMP.scala 361:36 362:17]
  wire  _GEN_3297 = cnt[6] ? _GEN_3280 : _GEN_3198; // @[NulCtrlMP.scala 708:22]
  wire  _GEN_3298 = cnt[6] ? _GEN_3281 : _GEN_3199; // @[NulCtrlMP.scala 708:22]
  wire  _GEN_3299 = cnt[6] ? _GEN_3282 : _GEN_3200; // @[NulCtrlMP.scala 708:22]
  wire  _GEN_3300 = cnt[6] ? _GEN_3283 : _GEN_3201; // @[NulCtrlMP.scala 708:22]
  wire [4:0] _GEN_3301 = cnt[6] ? _GEN_3284 : _GEN_3225; // @[NulCtrlMP.scala 708:22]
  wire [4:0] _GEN_3302 = cnt[6] ? _GEN_3285 : _GEN_3226; // @[NulCtrlMP.scala 708:22]
  wire [4:0] _GEN_3303 = cnt[6] ? _GEN_3286 : _GEN_3227; // @[NulCtrlMP.scala 708:22]
  wire [4:0] _GEN_3304 = cnt[6] ? _GEN_3287 : _GEN_3228; // @[NulCtrlMP.scala 708:22]
  wire [128:0] _GEN_3305 = cnt[6] ? _GEN_3288 : _GEN_3279; // @[NulCtrlMP.scala 708:22]
  wire  _GEN_3314 = _GEN_145 | _GEN_3221; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3315 = _GEN_146 | _GEN_3222; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3316 = _GEN_147 | _GEN_3223; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3317 = _GEN_148 | _GEN_3224; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_3318 = 2'h0 == opidx ? 5'h5 : _GEN_3301; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3319 = 2'h1 == opidx ? 5'h5 : _GEN_3302; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3320 = 2'h2 == opidx ? 5'h5 : _GEN_3303; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3321 = 2'h3 == opidx ? 5'h5 : _GEN_3304; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_3322 = 2'h0 == opidx ? regback_0 : _GEN_3229; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3323 = 2'h1 == opidx ? regback_0 : _GEN_3230; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3324 = 2'h2 == opidx ? regback_0 : _GEN_3231; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3325 = 2'h3 == opidx ? regback_0 : _GEN_3232; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_3326 = ~_GEN_1128 ? _cnt_T : _GEN_3305; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_3327 = cnt[7] ? _GEN_3314 : _GEN_3221; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3328 = cnt[7] ? _GEN_3315 : _GEN_3222; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3329 = cnt[7] ? _GEN_3316 : _GEN_3223; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3330 = cnt[7] ? _GEN_3317 : _GEN_3224; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3331 = cnt[7] ? _GEN_3318 : _GEN_3301; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3332 = cnt[7] ? _GEN_3319 : _GEN_3302; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3333 = cnt[7] ? _GEN_3320 : _GEN_3303; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3334 = cnt[7] ? _GEN_3321 : _GEN_3304; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3335 = cnt[7] ? _GEN_3322 : _GEN_3229; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3336 = cnt[7] ? _GEN_3323 : _GEN_3230; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3337 = cnt[7] ? _GEN_3324 : _GEN_3231; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3338 = cnt[7] ? _GEN_3325 : _GEN_3232; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3339 = cnt[7] ? _GEN_3326 : _GEN_3305; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3340 = _GEN_145 | _GEN_3327; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3341 = _GEN_146 | _GEN_3328; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3342 = _GEN_147 | _GEN_3329; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3343 = _GEN_148 | _GEN_3330; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_3344 = 2'h0 == opidx ? 5'h6 : _GEN_3331; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3345 = 2'h1 == opidx ? 5'h6 : _GEN_3332; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3346 = 2'h2 == opidx ? 5'h6 : _GEN_3333; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3347 = 2'h3 == opidx ? 5'h6 : _GEN_3334; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_3348 = 2'h0 == opidx ? regback_1 : _GEN_3335; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3349 = 2'h1 == opidx ? regback_1 : _GEN_3336; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3350 = 2'h2 == opidx ? regback_1 : _GEN_3337; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3351 = 2'h3 == opidx ? regback_1 : _GEN_3338; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_3352 = ~_GEN_1128 ? _cnt_T : _GEN_3339; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_3353 = cnt[8] ? _GEN_3340 : _GEN_3327; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3354 = cnt[8] ? _GEN_3341 : _GEN_3328; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3355 = cnt[8] ? _GEN_3342 : _GEN_3329; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3356 = cnt[8] ? _GEN_3343 : _GEN_3330; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3357 = cnt[8] ? _GEN_3344 : _GEN_3331; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3358 = cnt[8] ? _GEN_3345 : _GEN_3332; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3359 = cnt[8] ? _GEN_3346 : _GEN_3333; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3360 = cnt[8] ? _GEN_3347 : _GEN_3334; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3361 = cnt[8] ? _GEN_3348 : _GEN_3335; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3362 = cnt[8] ? _GEN_3349 : _GEN_3336; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3363 = cnt[8] ? _GEN_3350 : _GEN_3337; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3364 = cnt[8] ? _GEN_3351 : _GEN_3338; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3365 = cnt[8] ? _GEN_3352 : _GEN_3339; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3366 = cnt[9] ? 129'h1 : _GEN_3365; // @[NulCtrlMP.scala 710:22 711:17]
  wire [4:0] _GEN_3367 = cnt[9] ? 5'h5 : _GEN_3167; // @[NulCtrlMP.scala 710:22 712:19]
  wire  _GEN_3368 = state == 5'h10 ? _GEN_3297 : _GEN_3128; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3369 = state == 5'h10 ? _GEN_3298 : _GEN_3129; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3370 = state == 5'h10 ? _GEN_3299 : _GEN_3130; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3371 = state == 5'h10 ? _GEN_3300 : _GEN_3131; // @[NulCtrlMP.scala 702:33]
  wire [4:0] _GEN_3372 = state == 5'h10 ? _GEN_3357 : _GEN_3132; // @[NulCtrlMP.scala 702:33]
  wire [4:0] _GEN_3373 = state == 5'h10 ? _GEN_3358 : _GEN_3133; // @[NulCtrlMP.scala 702:33]
  wire [4:0] _GEN_3374 = state == 5'h10 ? _GEN_3359 : _GEN_3134; // @[NulCtrlMP.scala 702:33]
  wire [4:0] _GEN_3375 = state == 5'h10 ? _GEN_3360 : _GEN_3135; // @[NulCtrlMP.scala 702:33]
  wire [128:0] _GEN_3376 = state == 5'h10 ? _GEN_3366 : _GEN_3136; // @[NulCtrlMP.scala 702:33]
  wire [63:0] _GEN_3377 = state == 5'h10 ? _GEN_3187 : _GEN_3137; // @[NulCtrlMP.scala 702:33]
  wire [63:0] _GEN_3378 = state == 5'h10 ? _GEN_3207 : _GEN_3138; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3379 = state == 5'h10 ? _GEN_3353 : _GEN_3139; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3380 = state == 5'h10 ? _GEN_3354 : _GEN_3140; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3381 = state == 5'h10 ? _GEN_3355 : _GEN_3141; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3382 = state == 5'h10 ? _GEN_3356 : _GEN_3142; // @[NulCtrlMP.scala 702:33]
  wire [63:0] _GEN_3383 = state == 5'h10 ? _GEN_3361 : _GEN_3143; // @[NulCtrlMP.scala 702:33]
  wire [63:0] _GEN_3384 = state == 5'h10 ? _GEN_3362 : _GEN_3144; // @[NulCtrlMP.scala 702:33]
  wire [63:0] _GEN_3385 = state == 5'h10 ? _GEN_3363 : _GEN_3145; // @[NulCtrlMP.scala 702:33]
  wire [63:0] _GEN_3386 = state == 5'h10 ? _GEN_3364 : _GEN_3146; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3387 = state == 5'h10 ? _GEN_3261 : _GEN_3147; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3388 = state == 5'h10 ? _GEN_3262 : _GEN_3148; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3389 = state == 5'h10 ? _GEN_3263 : _GEN_3149; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3390 = state == 5'h10 ? _GEN_3264 : _GEN_3150; // @[NulCtrlMP.scala 702:33]
  wire [31:0] _GEN_3391 = state == 5'h10 ? _GEN_3265 : _GEN_3151; // @[NulCtrlMP.scala 702:33]
  wire [31:0] _GEN_3392 = state == 5'h10 ? _GEN_3266 : _GEN_3152; // @[NulCtrlMP.scala 702:33]
  wire [31:0] _GEN_3393 = state == 5'h10 ? _GEN_3267 : _GEN_3153; // @[NulCtrlMP.scala 702:33]
  wire [31:0] _GEN_3394 = state == 5'h10 ? _GEN_3268 : _GEN_3154; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3395 = state == 5'h10 ? _GEN_3275 : _GEN_3155; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3396 = state == 5'h10 ? _GEN_3276 : _GEN_3156; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3397 = state == 5'h10 ? _GEN_3277 : _GEN_3157; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3398 = state == 5'h10 ? _GEN_3278 : _GEN_3158; // @[NulCtrlMP.scala 702:33]
  wire [4:0] _GEN_3407 = state == 5'h10 ? _GEN_3367 : _GEN_3167; // @[NulCtrlMP.scala 702:33]
  wire  _GEN_3408 = _GEN_145 | _GEN_3368; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3409 = _GEN_146 | _GEN_3369; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3410 = _GEN_147 | _GEN_3370; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3411 = _GEN_148 | _GEN_3371; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_3412 = 2'h0 == opidx ? 5'h5 : _GEN_3372; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3413 = 2'h1 == opidx ? 5'h5 : _GEN_3373; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3414 = 2'h2 == opidx ? 5'h5 : _GEN_3374; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3415 = 2'h3 == opidx ? 5'h5 : _GEN_3375; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_3416 = _T_122 ? _cnt_T : _GEN_3376; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_3417 = _T_122 ? _GEN_1349 : _GEN_3377; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_3418 = cnt[0] ? _GEN_3408 : _GEN_3368; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3419 = cnt[0] ? _GEN_3409 : _GEN_3369; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3420 = cnt[0] ? _GEN_3410 : _GEN_3370; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3421 = cnt[0] ? _GEN_3411 : _GEN_3371; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3422 = cnt[0] ? _GEN_3412 : _GEN_3372; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3423 = cnt[0] ? _GEN_3413 : _GEN_3373; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3424 = cnt[0] ? _GEN_3414 : _GEN_3374; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3425 = cnt[0] ? _GEN_3415 : _GEN_3375; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_3426 = cnt[0] ? _GEN_3416 : _GEN_3376; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_3427 = cnt[0] ? _GEN_3417 : _GEN_3377; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3428 = _GEN_145 | _GEN_3418; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3429 = _GEN_146 | _GEN_3419; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3430 = _GEN_147 | _GEN_3420; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3431 = _GEN_148 | _GEN_3421; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_3432 = 2'h0 == opidx ? 5'h6 : _GEN_3422; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3433 = 2'h1 == opidx ? 5'h6 : _GEN_3423; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3434 = 2'h2 == opidx ? 5'h6 : _GEN_3424; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3435 = 2'h3 == opidx ? 5'h6 : _GEN_3425; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_3436 = _T_122 ? _cnt_T : _GEN_3426; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_3437 = _T_122 ? _GEN_1349 : _GEN_3378; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_3438 = cnt[1] ? _GEN_3428 : _GEN_3418; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3439 = cnt[1] ? _GEN_3429 : _GEN_3419; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3440 = cnt[1] ? _GEN_3430 : _GEN_3420; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3441 = cnt[1] ? _GEN_3431 : _GEN_3421; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3442 = cnt[1] ? _GEN_3432 : _GEN_3422; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3443 = cnt[1] ? _GEN_3433 : _GEN_3423; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3444 = cnt[1] ? _GEN_3434 : _GEN_3424; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3445 = cnt[1] ? _GEN_3435 : _GEN_3425; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_3446 = cnt[1] ? _GEN_3436 : _GEN_3426; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_3447 = cnt[1] ? _GEN_3437 : _GEN_3378; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3448 = _GEN_145 | _GEN_3379; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3449 = _GEN_146 | _GEN_3380; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3450 = _GEN_147 | _GEN_3381; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3451 = _GEN_148 | _GEN_3382; // @[NulCtrlMP.scala 377:{27,27}]
  wire [4:0] _GEN_3452 = 2'h0 == opidx ? 5'h5 : _GEN_3442; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3453 = 2'h1 == opidx ? 5'h5 : _GEN_3443; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3454 = 2'h2 == opidx ? 5'h5 : _GEN_3444; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3455 = 2'h3 == opidx ? 5'h5 : _GEN_3445; // @[NulCtrlMP.scala 378:{28,28}]
  wire [63:0] _GEN_3456 = 2'h0 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_3383; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3457 = 2'h1 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_3384; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3458 = 2'h2 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_3385; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3459 = 2'h3 == opidx ? _io_cpu_regacc_wdata_T_2 : _GEN_3386; // @[NulCtrlMP.scala 388:{30,30}]
  wire [128:0] _GEN_3460 = _T_122 ? _cnt_T : _GEN_3446; // @[NulCtrlMP.scala 389:36 390:17]
  wire  _GEN_3461 = cnt[2] ? _GEN_3448 : _GEN_3379; // @[NulCtrlMP.scala 718:22]
  wire  _GEN_3462 = cnt[2] ? _GEN_3449 : _GEN_3380; // @[NulCtrlMP.scala 718:22]
  wire  _GEN_3463 = cnt[2] ? _GEN_3450 : _GEN_3381; // @[NulCtrlMP.scala 718:22]
  wire  _GEN_3464 = cnt[2] ? _GEN_3451 : _GEN_3382; // @[NulCtrlMP.scala 718:22]
  wire [4:0] _GEN_3465 = cnt[2] ? _GEN_3452 : _GEN_3442; // @[NulCtrlMP.scala 718:22]
  wire [4:0] _GEN_3466 = cnt[2] ? _GEN_3453 : _GEN_3443; // @[NulCtrlMP.scala 718:22]
  wire [4:0] _GEN_3467 = cnt[2] ? _GEN_3454 : _GEN_3444; // @[NulCtrlMP.scala 718:22]
  wire [4:0] _GEN_3468 = cnt[2] ? _GEN_3455 : _GEN_3445; // @[NulCtrlMP.scala 718:22]
  wire [63:0] _GEN_3469 = cnt[2] ? _GEN_3456 : _GEN_3383; // @[NulCtrlMP.scala 718:22]
  wire [63:0] _GEN_3470 = cnt[2] ? _GEN_3457 : _GEN_3384; // @[NulCtrlMP.scala 718:22]
  wire [63:0] _GEN_3471 = cnt[2] ? _GEN_3458 : _GEN_3385; // @[NulCtrlMP.scala 718:22]
  wire [63:0] _GEN_3472 = cnt[2] ? _GEN_3459 : _GEN_3386; // @[NulCtrlMP.scala 718:22]
  wire [128:0] _GEN_3473 = cnt[2] ? _GEN_3460 : _GEN_3446; // @[NulCtrlMP.scala 718:22]
  wire  _GEN_3474 = _GEN_145 | _GEN_3461; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3475 = _GEN_146 | _GEN_3462; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3476 = _GEN_147 | _GEN_3463; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3477 = _GEN_148 | _GEN_3464; // @[NulCtrlMP.scala 377:{27,27}]
  wire [4:0] _GEN_3478 = 2'h0 == opidx ? 5'h6 : _GEN_3465; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3479 = 2'h1 == opidx ? 5'h6 : _GEN_3466; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3480 = 2'h2 == opidx ? 5'h6 : _GEN_3467; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3481 = 2'h3 == opidx ? 5'h6 : _GEN_3468; // @[NulCtrlMP.scala 378:{28,28}]
  wire [63:0] _io_cpu_regacc_wdata_T_5 = {oparg_15,oparg_14,oparg_13,oparg_12,oparg_11,oparg_10,oparg_9,oparg_8}; // @[NulCtrlMP.scala 388:53]
  wire [63:0] _GEN_3482 = 2'h0 == opidx ? _io_cpu_regacc_wdata_T_5 : _GEN_3469; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3483 = 2'h1 == opidx ? _io_cpu_regacc_wdata_T_5 : _GEN_3470; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3484 = 2'h2 == opidx ? _io_cpu_regacc_wdata_T_5 : _GEN_3471; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3485 = 2'h3 == opidx ? _io_cpu_regacc_wdata_T_5 : _GEN_3472; // @[NulCtrlMP.scala 388:{30,30}]
  wire [128:0] _GEN_3486 = _T_122 ? _cnt_T : _GEN_3473; // @[NulCtrlMP.scala 389:36 390:17]
  wire  _GEN_3487 = cnt[3] ? _GEN_3474 : _GEN_3461; // @[NulCtrlMP.scala 719:22]
  wire  _GEN_3488 = cnt[3] ? _GEN_3475 : _GEN_3462; // @[NulCtrlMP.scala 719:22]
  wire  _GEN_3489 = cnt[3] ? _GEN_3476 : _GEN_3463; // @[NulCtrlMP.scala 719:22]
  wire  _GEN_3490 = cnt[3] ? _GEN_3477 : _GEN_3464; // @[NulCtrlMP.scala 719:22]
  wire [4:0] _GEN_3491 = cnt[3] ? _GEN_3478 : _GEN_3465; // @[NulCtrlMP.scala 719:22]
  wire [4:0] _GEN_3492 = cnt[3] ? _GEN_3479 : _GEN_3466; // @[NulCtrlMP.scala 719:22]
  wire [4:0] _GEN_3493 = cnt[3] ? _GEN_3480 : _GEN_3467; // @[NulCtrlMP.scala 719:22]
  wire [4:0] _GEN_3494 = cnt[3] ? _GEN_3481 : _GEN_3468; // @[NulCtrlMP.scala 719:22]
  wire [63:0] _GEN_3495 = cnt[3] ? _GEN_3482 : _GEN_3469; // @[NulCtrlMP.scala 719:22]
  wire [63:0] _GEN_3496 = cnt[3] ? _GEN_3483 : _GEN_3470; // @[NulCtrlMP.scala 719:22]
  wire [63:0] _GEN_3497 = cnt[3] ? _GEN_3484 : _GEN_3471; // @[NulCtrlMP.scala 719:22]
  wire [63:0] _GEN_3498 = cnt[3] ? _GEN_3485 : _GEN_3472; // @[NulCtrlMP.scala 719:22]
  wire [128:0] _GEN_3499 = cnt[3] ? _GEN_3486 : _GEN_3473; // @[NulCtrlMP.scala 719:22]
  wire  _GEN_3500 = _GEN_145 | _GEN_3387; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3501 = _GEN_146 | _GEN_3388; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3502 = _GEN_147 | _GEN_3389; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3503 = _GEN_148 | _GEN_3390; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3504 = 2'h0 == opidx ? 32'h62b023 : _GEN_3391; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3505 = 2'h1 == opidx ? 32'h62b023 : _GEN_3392; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3506 = 2'h2 == opidx ? 32'h62b023 : _GEN_3393; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3507 = 2'h3 == opidx ? 32'h62b023 : _GEN_3394; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3508 = _GEN_1180 ? _cnt_T : _GEN_3499; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3509 = cnt[4] ? _GEN_3500 : _GEN_3387; // @[NulCtrlMP.scala 720:22]
  wire  _GEN_3510 = cnt[4] ? _GEN_3501 : _GEN_3388; // @[NulCtrlMP.scala 720:22]
  wire  _GEN_3511 = cnt[4] ? _GEN_3502 : _GEN_3389; // @[NulCtrlMP.scala 720:22]
  wire  _GEN_3512 = cnt[4] ? _GEN_3503 : _GEN_3390; // @[NulCtrlMP.scala 720:22]
  wire [31:0] _GEN_3513 = cnt[4] ? _GEN_3504 : _GEN_3391; // @[NulCtrlMP.scala 720:22]
  wire [31:0] _GEN_3514 = cnt[4] ? _GEN_3505 : _GEN_3392; // @[NulCtrlMP.scala 720:22]
  wire [31:0] _GEN_3515 = cnt[4] ? _GEN_3506 : _GEN_3393; // @[NulCtrlMP.scala 720:22]
  wire [31:0] _GEN_3516 = cnt[4] ? _GEN_3507 : _GEN_3394; // @[NulCtrlMP.scala 720:22]
  wire [128:0] _GEN_3517 = cnt[4] ? _GEN_3508 : _GEN_3499; // @[NulCtrlMP.scala 720:22]
  wire  _GEN_3518 = _GEN_145 | _GEN_3509; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3519 = _GEN_146 | _GEN_3510; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3520 = _GEN_147 | _GEN_3511; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3521 = _GEN_148 | _GEN_3512; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3522 = 2'h0 == opidx ? 32'h330000f : _GEN_3513; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3523 = 2'h1 == opidx ? 32'h330000f : _GEN_3514; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3524 = 2'h2 == opidx ? 32'h330000f : _GEN_3515; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3525 = 2'h3 == opidx ? 32'h330000f : _GEN_3516; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3526 = _GEN_1180 ? _cnt_T : _GEN_3517; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3527 = cnt[5] ? _GEN_3518 : _GEN_3509; // @[NulCtrlMP.scala 721:22]
  wire  _GEN_3528 = cnt[5] ? _GEN_3519 : _GEN_3510; // @[NulCtrlMP.scala 721:22]
  wire  _GEN_3529 = cnt[5] ? _GEN_3520 : _GEN_3511; // @[NulCtrlMP.scala 721:22]
  wire  _GEN_3530 = cnt[5] ? _GEN_3521 : _GEN_3512; // @[NulCtrlMP.scala 721:22]
  wire [31:0] _GEN_3531 = cnt[5] ? _GEN_3522 : _GEN_3513; // @[NulCtrlMP.scala 721:22]
  wire [31:0] _GEN_3532 = cnt[5] ? _GEN_3523 : _GEN_3514; // @[NulCtrlMP.scala 721:22]
  wire [31:0] _GEN_3533 = cnt[5] ? _GEN_3524 : _GEN_3515; // @[NulCtrlMP.scala 721:22]
  wire [31:0] _GEN_3534 = cnt[5] ? _GEN_3525 : _GEN_3516; // @[NulCtrlMP.scala 721:22]
  wire [128:0] _GEN_3535 = cnt[5] ? _GEN_3526 : _GEN_3517; // @[NulCtrlMP.scala 721:22]
  wire  _GEN_3536 = _GEN_145 | _GEN_3395; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3537 = _GEN_146 | _GEN_3396; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3538 = _GEN_147 | _GEN_3397; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3539 = _GEN_148 | _GEN_3398; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_3540 = ~_GEN_1252 ? _cnt_T : _GEN_3535; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_3541 = cnt[6] ? _GEN_3536 : _GEN_3395; // @[NulCtrlMP.scala 722:22]
  wire  _GEN_3542 = cnt[6] ? _GEN_3537 : _GEN_3396; // @[NulCtrlMP.scala 722:22]
  wire  _GEN_3543 = cnt[6] ? _GEN_3538 : _GEN_3397; // @[NulCtrlMP.scala 722:22]
  wire  _GEN_3544 = cnt[6] ? _GEN_3539 : _GEN_3398; // @[NulCtrlMP.scala 722:22]
  wire [128:0] _GEN_3545 = cnt[6] ? _GEN_3540 : _GEN_3535; // @[NulCtrlMP.scala 722:22]
  wire  _GEN_3546 = _GEN_145 | _GEN_3487; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3547 = _GEN_146 | _GEN_3488; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3548 = _GEN_147 | _GEN_3489; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3549 = _GEN_148 | _GEN_3490; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_3550 = 2'h0 == opidx ? 5'h5 : _GEN_3491; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3551 = 2'h1 == opidx ? 5'h5 : _GEN_3492; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3552 = 2'h2 == opidx ? 5'h5 : _GEN_3493; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3553 = 2'h3 == opidx ? 5'h5 : _GEN_3494; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_3554 = 2'h0 == opidx ? regback_0 : _GEN_3495; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3555 = 2'h1 == opidx ? regback_0 : _GEN_3496; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3556 = 2'h2 == opidx ? regback_0 : _GEN_3497; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3557 = 2'h3 == opidx ? regback_0 : _GEN_3498; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_3558 = ~_GEN_1128 ? _cnt_T : _GEN_3545; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_3559 = cnt[7] ? _GEN_3546 : _GEN_3487; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3560 = cnt[7] ? _GEN_3547 : _GEN_3488; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3561 = cnt[7] ? _GEN_3548 : _GEN_3489; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3562 = cnt[7] ? _GEN_3549 : _GEN_3490; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3563 = cnt[7] ? _GEN_3550 : _GEN_3491; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3564 = cnt[7] ? _GEN_3551 : _GEN_3492; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3565 = cnt[7] ? _GEN_3552 : _GEN_3493; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3566 = cnt[7] ? _GEN_3553 : _GEN_3494; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3567 = cnt[7] ? _GEN_3554 : _GEN_3495; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3568 = cnt[7] ? _GEN_3555 : _GEN_3496; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3569 = cnt[7] ? _GEN_3556 : _GEN_3497; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3570 = cnt[7] ? _GEN_3557 : _GEN_3498; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3571 = cnt[7] ? _GEN_3558 : _GEN_3545; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3572 = _GEN_145 | _GEN_3559; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3573 = _GEN_146 | _GEN_3560; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3574 = _GEN_147 | _GEN_3561; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3575 = _GEN_148 | _GEN_3562; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_3576 = 2'h0 == opidx ? 5'h6 : _GEN_3563; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3577 = 2'h1 == opidx ? 5'h6 : _GEN_3564; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3578 = 2'h2 == opidx ? 5'h6 : _GEN_3565; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3579 = 2'h3 == opidx ? 5'h6 : _GEN_3566; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_3580 = 2'h0 == opidx ? regback_1 : _GEN_3567; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3581 = 2'h1 == opidx ? regback_1 : _GEN_3568; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3582 = 2'h2 == opidx ? regback_1 : _GEN_3569; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3583 = 2'h3 == opidx ? regback_1 : _GEN_3570; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_3584 = ~_GEN_1128 ? _cnt_T : _GEN_3571; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_3585 = cnt[8] ? _GEN_3572 : _GEN_3559; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3586 = cnt[8] ? _GEN_3573 : _GEN_3560; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3587 = cnt[8] ? _GEN_3574 : _GEN_3561; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3588 = cnt[8] ? _GEN_3575 : _GEN_3562; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3589 = cnt[8] ? _GEN_3576 : _GEN_3563; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3590 = cnt[8] ? _GEN_3577 : _GEN_3564; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3591 = cnt[8] ? _GEN_3578 : _GEN_3565; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3592 = cnt[8] ? _GEN_3579 : _GEN_3566; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3593 = cnt[8] ? _GEN_3580 : _GEN_3567; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3594 = cnt[8] ? _GEN_3581 : _GEN_3568; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3595 = cnt[8] ? _GEN_3582 : _GEN_3569; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3596 = cnt[8] ? _GEN_3583 : _GEN_3570; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3597 = cnt[8] ? _GEN_3584 : _GEN_3571; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3598 = cnt[9] ? 129'h1 : _GEN_3597; // @[NulCtrlMP.scala 724:22 725:17]
  wire [4:0] _GEN_3599 = cnt[9] ? 5'h5 : _GEN_3407; // @[NulCtrlMP.scala 724:22 726:19]
  wire  _GEN_3600 = state == 5'h11 ? _GEN_3438 : _GEN_3368; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3601 = state == 5'h11 ? _GEN_3439 : _GEN_3369; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3602 = state == 5'h11 ? _GEN_3440 : _GEN_3370; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3603 = state == 5'h11 ? _GEN_3441 : _GEN_3371; // @[NulCtrlMP.scala 716:33]
  wire [4:0] _GEN_3604 = state == 5'h11 ? _GEN_3589 : _GEN_3372; // @[NulCtrlMP.scala 716:33]
  wire [4:0] _GEN_3605 = state == 5'h11 ? _GEN_3590 : _GEN_3373; // @[NulCtrlMP.scala 716:33]
  wire [4:0] _GEN_3606 = state == 5'h11 ? _GEN_3591 : _GEN_3374; // @[NulCtrlMP.scala 716:33]
  wire [4:0] _GEN_3607 = state == 5'h11 ? _GEN_3592 : _GEN_3375; // @[NulCtrlMP.scala 716:33]
  wire [128:0] _GEN_3608 = state == 5'h11 ? _GEN_3598 : _GEN_3376; // @[NulCtrlMP.scala 716:33]
  wire [63:0] _GEN_3609 = state == 5'h11 ? _GEN_3427 : _GEN_3377; // @[NulCtrlMP.scala 716:33]
  wire [63:0] _GEN_3610 = state == 5'h11 ? _GEN_3447 : _GEN_3378; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3611 = state == 5'h11 ? _GEN_3585 : _GEN_3379; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3612 = state == 5'h11 ? _GEN_3586 : _GEN_3380; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3613 = state == 5'h11 ? _GEN_3587 : _GEN_3381; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3614 = state == 5'h11 ? _GEN_3588 : _GEN_3382; // @[NulCtrlMP.scala 716:33]
  wire [63:0] _GEN_3615 = state == 5'h11 ? _GEN_3593 : _GEN_3383; // @[NulCtrlMP.scala 716:33]
  wire [63:0] _GEN_3616 = state == 5'h11 ? _GEN_3594 : _GEN_3384; // @[NulCtrlMP.scala 716:33]
  wire [63:0] _GEN_3617 = state == 5'h11 ? _GEN_3595 : _GEN_3385; // @[NulCtrlMP.scala 716:33]
  wire [63:0] _GEN_3618 = state == 5'h11 ? _GEN_3596 : _GEN_3386; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3619 = state == 5'h11 ? _GEN_3527 : _GEN_3387; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3620 = state == 5'h11 ? _GEN_3528 : _GEN_3388; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3621 = state == 5'h11 ? _GEN_3529 : _GEN_3389; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3622 = state == 5'h11 ? _GEN_3530 : _GEN_3390; // @[NulCtrlMP.scala 716:33]
  wire [31:0] _GEN_3623 = state == 5'h11 ? _GEN_3531 : _GEN_3391; // @[NulCtrlMP.scala 716:33]
  wire [31:0] _GEN_3624 = state == 5'h11 ? _GEN_3532 : _GEN_3392; // @[NulCtrlMP.scala 716:33]
  wire [31:0] _GEN_3625 = state == 5'h11 ? _GEN_3533 : _GEN_3393; // @[NulCtrlMP.scala 716:33]
  wire [31:0] _GEN_3626 = state == 5'h11 ? _GEN_3534 : _GEN_3394; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3627 = state == 5'h11 ? _GEN_3541 : _GEN_3395; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3628 = state == 5'h11 ? _GEN_3542 : _GEN_3396; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3629 = state == 5'h11 ? _GEN_3543 : _GEN_3397; // @[NulCtrlMP.scala 716:33]
  wire  _GEN_3630 = state == 5'h11 ? _GEN_3544 : _GEN_3398; // @[NulCtrlMP.scala 716:33]
  wire [4:0] _GEN_3631 = state == 5'h11 ? _GEN_3599 : _GEN_3407; // @[NulCtrlMP.scala 716:33]
  wire [63:0] pg_base_addr2 = {12'h0,oparg_6,oparg_5,oparg_4,oparg_3,oparg_2,12'h0}; // @[Cat.scala 31:58]
  wire [63:0] pg_base_addr7 = {12'h0,oparg_11,oparg_10,oparg_9,oparg_8,oparg_7,12'h0}; // @[Cat.scala 31:58]
  reg [7:0] pg_loop_cnt; // @[NulCtrlMP.scala 742:30]
  wire  _GEN_3632 = _GEN_145 | _GEN_3600; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3633 = _GEN_146 | _GEN_3601; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3634 = _GEN_147 | _GEN_3602; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3635 = _GEN_148 | _GEN_3603; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_3636 = 2'h0 == opidx ? 5'h5 : _GEN_3604; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3637 = 2'h1 == opidx ? 5'h5 : _GEN_3605; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3638 = 2'h2 == opidx ? 5'h5 : _GEN_3606; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3639 = 2'h3 == opidx ? 5'h5 : _GEN_3607; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_3640 = _T_122 ? _cnt_T : _GEN_3608; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_3641 = _T_122 ? _GEN_1349 : _GEN_3609; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_3642 = cnt[0] ? _GEN_3632 : _GEN_3600; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3643 = cnt[0] ? _GEN_3633 : _GEN_3601; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3644 = cnt[0] ? _GEN_3634 : _GEN_3602; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3645 = cnt[0] ? _GEN_3635 : _GEN_3603; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3646 = cnt[0] ? _GEN_3636 : _GEN_3604; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3647 = cnt[0] ? _GEN_3637 : _GEN_3605; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3648 = cnt[0] ? _GEN_3638 : _GEN_3606; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3649 = cnt[0] ? _GEN_3639 : _GEN_3607; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_3650 = cnt[0] ? _GEN_3640 : _GEN_3608; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_3651 = cnt[0] ? _GEN_3641 : _GEN_3609; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3652 = _GEN_145 | _GEN_3642; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3653 = _GEN_146 | _GEN_3643; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3654 = _GEN_147 | _GEN_3644; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_3655 = _GEN_148 | _GEN_3645; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_3656 = 2'h0 == opidx ? 5'h6 : _GEN_3646; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3657 = 2'h1 == opidx ? 5'h6 : _GEN_3647; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3658 = 2'h2 == opidx ? 5'h6 : _GEN_3648; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_3659 = 2'h3 == opidx ? 5'h6 : _GEN_3649; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_3660 = _T_122 ? _cnt_T : _GEN_3650; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_3661 = _T_122 ? _GEN_1349 : _GEN_3610; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_3662 = cnt[1] ? _GEN_3652 : _GEN_3642; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3663 = cnt[1] ? _GEN_3653 : _GEN_3643; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3664 = cnt[1] ? _GEN_3654 : _GEN_3644; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3665 = cnt[1] ? _GEN_3655 : _GEN_3645; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3666 = cnt[1] ? _GEN_3656 : _GEN_3646; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3667 = cnt[1] ? _GEN_3657 : _GEN_3647; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3668 = cnt[1] ? _GEN_3658 : _GEN_3648; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_3669 = cnt[1] ? _GEN_3659 : _GEN_3649; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_3670 = cnt[1] ? _GEN_3660 : _GEN_3650; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_3671 = cnt[1] ? _GEN_3661 : _GEN_3610; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_3672 = _GEN_145 | _GEN_3611; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3673 = _GEN_146 | _GEN_3612; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3674 = _GEN_147 | _GEN_3613; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3675 = _GEN_148 | _GEN_3614; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_3676 = 2'h0 == opidx ? 5'h5 : _GEN_3666; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3677 = 2'h1 == opidx ? 5'h5 : _GEN_3667; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3678 = 2'h2 == opidx ? 5'h5 : _GEN_3668; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3679 = 2'h3 == opidx ? 5'h5 : _GEN_3669; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_3680 = 2'h0 == opidx ? pg_base_addr2 : _GEN_3615; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3681 = 2'h1 == opidx ? pg_base_addr2 : _GEN_3616; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3682 = 2'h2 == opidx ? pg_base_addr2 : _GEN_3617; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3683 = 2'h3 == opidx ? pg_base_addr2 : _GEN_3618; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_3684 = ~_GEN_1128 ? _cnt_T : _GEN_3670; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_3685 = cnt[2] ? _GEN_3672 : _GEN_3611; // @[NulCtrlMP.scala 747:22]
  wire  _GEN_3686 = cnt[2] ? _GEN_3673 : _GEN_3612; // @[NulCtrlMP.scala 747:22]
  wire  _GEN_3687 = cnt[2] ? _GEN_3674 : _GEN_3613; // @[NulCtrlMP.scala 747:22]
  wire  _GEN_3688 = cnt[2] ? _GEN_3675 : _GEN_3614; // @[NulCtrlMP.scala 747:22]
  wire [4:0] _GEN_3689 = cnt[2] ? _GEN_3676 : _GEN_3666; // @[NulCtrlMP.scala 747:22]
  wire [4:0] _GEN_3690 = cnt[2] ? _GEN_3677 : _GEN_3667; // @[NulCtrlMP.scala 747:22]
  wire [4:0] _GEN_3691 = cnt[2] ? _GEN_3678 : _GEN_3668; // @[NulCtrlMP.scala 747:22]
  wire [4:0] _GEN_3692 = cnt[2] ? _GEN_3679 : _GEN_3669; // @[NulCtrlMP.scala 747:22]
  wire [63:0] _GEN_3693 = cnt[2] ? _GEN_3680 : _GEN_3615; // @[NulCtrlMP.scala 747:22]
  wire [63:0] _GEN_3694 = cnt[2] ? _GEN_3681 : _GEN_3616; // @[NulCtrlMP.scala 747:22]
  wire [63:0] _GEN_3695 = cnt[2] ? _GEN_3682 : _GEN_3617; // @[NulCtrlMP.scala 747:22]
  wire [63:0] _GEN_3696 = cnt[2] ? _GEN_3683 : _GEN_3618; // @[NulCtrlMP.scala 747:22]
  wire [128:0] _GEN_3697 = cnt[2] ? _GEN_3684 : _GEN_3670; // @[NulCtrlMP.scala 747:22]
  wire  _GEN_3698 = _GEN_145 | _GEN_3685; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3699 = _GEN_146 | _GEN_3686; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3700 = _GEN_147 | _GEN_3687; // @[NulCtrlMP.scala 377:{27,27}]
  wire  _GEN_3701 = _GEN_148 | _GEN_3688; // @[NulCtrlMP.scala 377:{27,27}]
  wire [4:0] _GEN_3702 = 2'h0 == opidx ? 5'h6 : _GEN_3689; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3703 = 2'h1 == opidx ? 5'h6 : _GEN_3690; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3704 = 2'h2 == opidx ? 5'h6 : _GEN_3691; // @[NulCtrlMP.scala 378:{28,28}]
  wire [4:0] _GEN_3705 = 2'h3 == opidx ? 5'h6 : _GEN_3692; // @[NulCtrlMP.scala 378:{28,28}]
  wire [63:0] _io_cpu_regacc_wdata_T_6 = {oparg_14,oparg_13,oparg_12,oparg_11,oparg_10,oparg_9,oparg_8,oparg_7}; // @[NulCtrlMP.scala 388:53]
  wire [63:0] _GEN_3706 = 2'h0 == opidx ? _io_cpu_regacc_wdata_T_6 : _GEN_3693; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3707 = 2'h1 == opidx ? _io_cpu_regacc_wdata_T_6 : _GEN_3694; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3708 = 2'h2 == opidx ? _io_cpu_regacc_wdata_T_6 : _GEN_3695; // @[NulCtrlMP.scala 388:{30,30}]
  wire [63:0] _GEN_3709 = 2'h3 == opidx ? _io_cpu_regacc_wdata_T_6 : _GEN_3696; // @[NulCtrlMP.scala 388:{30,30}]
  wire [128:0] _GEN_3710 = _T_122 ? _cnt_T : _GEN_3697; // @[NulCtrlMP.scala 389:36 390:17]
  wire  _GEN_3711 = cnt[3] ? _GEN_3698 : _GEN_3685; // @[NulCtrlMP.scala 748:22]
  wire  _GEN_3712 = cnt[3] ? _GEN_3699 : _GEN_3686; // @[NulCtrlMP.scala 748:22]
  wire  _GEN_3713 = cnt[3] ? _GEN_3700 : _GEN_3687; // @[NulCtrlMP.scala 748:22]
  wire  _GEN_3714 = cnt[3] ? _GEN_3701 : _GEN_3688; // @[NulCtrlMP.scala 748:22]
  wire [4:0] _GEN_3715 = cnt[3] ? _GEN_3702 : _GEN_3689; // @[NulCtrlMP.scala 748:22]
  wire [4:0] _GEN_3716 = cnt[3] ? _GEN_3703 : _GEN_3690; // @[NulCtrlMP.scala 748:22]
  wire [4:0] _GEN_3717 = cnt[3] ? _GEN_3704 : _GEN_3691; // @[NulCtrlMP.scala 748:22]
  wire [4:0] _GEN_3718 = cnt[3] ? _GEN_3705 : _GEN_3692; // @[NulCtrlMP.scala 748:22]
  wire [63:0] _GEN_3719 = cnt[3] ? _GEN_3706 : _GEN_3693; // @[NulCtrlMP.scala 748:22]
  wire [63:0] _GEN_3720 = cnt[3] ? _GEN_3707 : _GEN_3694; // @[NulCtrlMP.scala 748:22]
  wire [63:0] _GEN_3721 = cnt[3] ? _GEN_3708 : _GEN_3695; // @[NulCtrlMP.scala 748:22]
  wire [63:0] _GEN_3722 = cnt[3] ? _GEN_3709 : _GEN_3696; // @[NulCtrlMP.scala 748:22]
  wire [128:0] _GEN_3723 = cnt[3] ? _GEN_3710 : _GEN_3697; // @[NulCtrlMP.scala 748:22]
  wire  _GEN_3724 = _GEN_145 | _GEN_3619; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3725 = _GEN_146 | _GEN_3620; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3726 = _GEN_147 | _GEN_3621; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3727 = _GEN_148 | _GEN_3622; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3728 = 2'h0 == opidx ? 32'h62b023 : _GEN_3623; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3729 = 2'h1 == opidx ? 32'h62b023 : _GEN_3624; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3730 = 2'h2 == opidx ? 32'h62b023 : _GEN_3625; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3731 = 2'h3 == opidx ? 32'h62b023 : _GEN_3626; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3732 = _GEN_1180 ? _cnt_T : _GEN_3723; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3733 = cnt[4] ? _GEN_3724 : _GEN_3619; // @[NulCtrlMP.scala 749:22]
  wire  _GEN_3734 = cnt[4] ? _GEN_3725 : _GEN_3620; // @[NulCtrlMP.scala 749:22]
  wire  _GEN_3735 = cnt[4] ? _GEN_3726 : _GEN_3621; // @[NulCtrlMP.scala 749:22]
  wire  _GEN_3736 = cnt[4] ? _GEN_3727 : _GEN_3622; // @[NulCtrlMP.scala 749:22]
  wire [31:0] _GEN_3737 = cnt[4] ? _GEN_3728 : _GEN_3623; // @[NulCtrlMP.scala 749:22]
  wire [31:0] _GEN_3738 = cnt[4] ? _GEN_3729 : _GEN_3624; // @[NulCtrlMP.scala 749:22]
  wire [31:0] _GEN_3739 = cnt[4] ? _GEN_3730 : _GEN_3625; // @[NulCtrlMP.scala 749:22]
  wire [31:0] _GEN_3740 = cnt[4] ? _GEN_3731 : _GEN_3626; // @[NulCtrlMP.scala 749:22]
  wire [128:0] _GEN_3741 = cnt[4] ? _GEN_3732 : _GEN_3723; // @[NulCtrlMP.scala 749:22]
  wire  _GEN_3742 = _GEN_145 | _GEN_3733; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3743 = _GEN_146 | _GEN_3734; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3744 = _GEN_147 | _GEN_3735; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3745 = _GEN_148 | _GEN_3736; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3746 = 2'h0 == opidx ? 32'h62b423 : _GEN_3737; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3747 = 2'h1 == opidx ? 32'h62b423 : _GEN_3738; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3748 = 2'h2 == opidx ? 32'h62b423 : _GEN_3739; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3749 = 2'h3 == opidx ? 32'h62b423 : _GEN_3740; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3750 = _GEN_1180 ? _cnt_T : _GEN_3741; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3751 = cnt[5] ? _GEN_3742 : _GEN_3733; // @[NulCtrlMP.scala 750:22]
  wire  _GEN_3752 = cnt[5] ? _GEN_3743 : _GEN_3734; // @[NulCtrlMP.scala 750:22]
  wire  _GEN_3753 = cnt[5] ? _GEN_3744 : _GEN_3735; // @[NulCtrlMP.scala 750:22]
  wire  _GEN_3754 = cnt[5] ? _GEN_3745 : _GEN_3736; // @[NulCtrlMP.scala 750:22]
  wire [31:0] _GEN_3755 = cnt[5] ? _GEN_3746 : _GEN_3737; // @[NulCtrlMP.scala 750:22]
  wire [31:0] _GEN_3756 = cnt[5] ? _GEN_3747 : _GEN_3738; // @[NulCtrlMP.scala 750:22]
  wire [31:0] _GEN_3757 = cnt[5] ? _GEN_3748 : _GEN_3739; // @[NulCtrlMP.scala 750:22]
  wire [31:0] _GEN_3758 = cnt[5] ? _GEN_3749 : _GEN_3740; // @[NulCtrlMP.scala 750:22]
  wire [128:0] _GEN_3759 = cnt[5] ? _GEN_3750 : _GEN_3741; // @[NulCtrlMP.scala 750:22]
  wire  _GEN_3760 = _GEN_145 | _GEN_3751; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3761 = _GEN_146 | _GEN_3752; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3762 = _GEN_147 | _GEN_3753; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3763 = _GEN_148 | _GEN_3754; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3764 = 2'h0 == opidx ? 32'h62b823 : _GEN_3755; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3765 = 2'h1 == opidx ? 32'h62b823 : _GEN_3756; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3766 = 2'h2 == opidx ? 32'h62b823 : _GEN_3757; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3767 = 2'h3 == opidx ? 32'h62b823 : _GEN_3758; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3768 = _GEN_1180 ? _cnt_T : _GEN_3759; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3769 = cnt[6] ? _GEN_3760 : _GEN_3751; // @[NulCtrlMP.scala 751:22]
  wire  _GEN_3770 = cnt[6] ? _GEN_3761 : _GEN_3752; // @[NulCtrlMP.scala 751:22]
  wire  _GEN_3771 = cnt[6] ? _GEN_3762 : _GEN_3753; // @[NulCtrlMP.scala 751:22]
  wire  _GEN_3772 = cnt[6] ? _GEN_3763 : _GEN_3754; // @[NulCtrlMP.scala 751:22]
  wire [31:0] _GEN_3773 = cnt[6] ? _GEN_3764 : _GEN_3755; // @[NulCtrlMP.scala 751:22]
  wire [31:0] _GEN_3774 = cnt[6] ? _GEN_3765 : _GEN_3756; // @[NulCtrlMP.scala 751:22]
  wire [31:0] _GEN_3775 = cnt[6] ? _GEN_3766 : _GEN_3757; // @[NulCtrlMP.scala 751:22]
  wire [31:0] _GEN_3776 = cnt[6] ? _GEN_3767 : _GEN_3758; // @[NulCtrlMP.scala 751:22]
  wire [128:0] _GEN_3777 = cnt[6] ? _GEN_3768 : _GEN_3759; // @[NulCtrlMP.scala 751:22]
  wire  _GEN_3778 = _GEN_145 | _GEN_3769; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3779 = _GEN_146 | _GEN_3770; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3780 = _GEN_147 | _GEN_3771; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3781 = _GEN_148 | _GEN_3772; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3782 = 2'h0 == opidx ? 32'h62bc23 : _GEN_3773; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3783 = 2'h1 == opidx ? 32'h62bc23 : _GEN_3774; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3784 = 2'h2 == opidx ? 32'h62bc23 : _GEN_3775; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3785 = 2'h3 == opidx ? 32'h62bc23 : _GEN_3776; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3786 = _GEN_1180 ? _cnt_T : _GEN_3777; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3787 = cnt[7] ? _GEN_3778 : _GEN_3769; // @[NulCtrlMP.scala 752:22]
  wire  _GEN_3788 = cnt[7] ? _GEN_3779 : _GEN_3770; // @[NulCtrlMP.scala 752:22]
  wire  _GEN_3789 = cnt[7] ? _GEN_3780 : _GEN_3771; // @[NulCtrlMP.scala 752:22]
  wire  _GEN_3790 = cnt[7] ? _GEN_3781 : _GEN_3772; // @[NulCtrlMP.scala 752:22]
  wire [31:0] _GEN_3791 = cnt[7] ? _GEN_3782 : _GEN_3773; // @[NulCtrlMP.scala 752:22]
  wire [31:0] _GEN_3792 = cnt[7] ? _GEN_3783 : _GEN_3774; // @[NulCtrlMP.scala 752:22]
  wire [31:0] _GEN_3793 = cnt[7] ? _GEN_3784 : _GEN_3775; // @[NulCtrlMP.scala 752:22]
  wire [31:0] _GEN_3794 = cnt[7] ? _GEN_3785 : _GEN_3776; // @[NulCtrlMP.scala 752:22]
  wire [128:0] _GEN_3795 = cnt[7] ? _GEN_3786 : _GEN_3777; // @[NulCtrlMP.scala 752:22]
  wire  _GEN_3796 = _GEN_145 | _GEN_3787; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3797 = _GEN_146 | _GEN_3788; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3798 = _GEN_147 | _GEN_3789; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3799 = _GEN_148 | _GEN_3790; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3800 = 2'h0 == opidx ? 32'h262b023 : _GEN_3791; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3801 = 2'h1 == opidx ? 32'h262b023 : _GEN_3792; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3802 = 2'h2 == opidx ? 32'h262b023 : _GEN_3793; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3803 = 2'h3 == opidx ? 32'h262b023 : _GEN_3794; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3804 = _GEN_1180 ? _cnt_T : _GEN_3795; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3805 = cnt[8] ? _GEN_3796 : _GEN_3787; // @[NulCtrlMP.scala 753:22]
  wire  _GEN_3806 = cnt[8] ? _GEN_3797 : _GEN_3788; // @[NulCtrlMP.scala 753:22]
  wire  _GEN_3807 = cnt[8] ? _GEN_3798 : _GEN_3789; // @[NulCtrlMP.scala 753:22]
  wire  _GEN_3808 = cnt[8] ? _GEN_3799 : _GEN_3790; // @[NulCtrlMP.scala 753:22]
  wire [31:0] _GEN_3809 = cnt[8] ? _GEN_3800 : _GEN_3791; // @[NulCtrlMP.scala 753:22]
  wire [31:0] _GEN_3810 = cnt[8] ? _GEN_3801 : _GEN_3792; // @[NulCtrlMP.scala 753:22]
  wire [31:0] _GEN_3811 = cnt[8] ? _GEN_3802 : _GEN_3793; // @[NulCtrlMP.scala 753:22]
  wire [31:0] _GEN_3812 = cnt[8] ? _GEN_3803 : _GEN_3794; // @[NulCtrlMP.scala 753:22]
  wire [128:0] _GEN_3813 = cnt[8] ? _GEN_3804 : _GEN_3795; // @[NulCtrlMP.scala 753:22]
  wire  _GEN_3814 = _GEN_145 | _GEN_3805; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3815 = _GEN_146 | _GEN_3806; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3816 = _GEN_147 | _GEN_3807; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3817 = _GEN_148 | _GEN_3808; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3818 = 2'h0 == opidx ? 32'h262b423 : _GEN_3809; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3819 = 2'h1 == opidx ? 32'h262b423 : _GEN_3810; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3820 = 2'h2 == opidx ? 32'h262b423 : _GEN_3811; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3821 = 2'h3 == opidx ? 32'h262b423 : _GEN_3812; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3822 = _GEN_1180 ? _cnt_T : _GEN_3813; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3823 = cnt[9] ? _GEN_3814 : _GEN_3805; // @[NulCtrlMP.scala 754:22]
  wire  _GEN_3824 = cnt[9] ? _GEN_3815 : _GEN_3806; // @[NulCtrlMP.scala 754:22]
  wire  _GEN_3825 = cnt[9] ? _GEN_3816 : _GEN_3807; // @[NulCtrlMP.scala 754:22]
  wire  _GEN_3826 = cnt[9] ? _GEN_3817 : _GEN_3808; // @[NulCtrlMP.scala 754:22]
  wire [31:0] _GEN_3827 = cnt[9] ? _GEN_3818 : _GEN_3809; // @[NulCtrlMP.scala 754:22]
  wire [31:0] _GEN_3828 = cnt[9] ? _GEN_3819 : _GEN_3810; // @[NulCtrlMP.scala 754:22]
  wire [31:0] _GEN_3829 = cnt[9] ? _GEN_3820 : _GEN_3811; // @[NulCtrlMP.scala 754:22]
  wire [31:0] _GEN_3830 = cnt[9] ? _GEN_3821 : _GEN_3812; // @[NulCtrlMP.scala 754:22]
  wire [128:0] _GEN_3831 = cnt[9] ? _GEN_3822 : _GEN_3813; // @[NulCtrlMP.scala 754:22]
  wire  _GEN_3832 = _GEN_145 | _GEN_3823; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3833 = _GEN_146 | _GEN_3824; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3834 = _GEN_147 | _GEN_3825; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3835 = _GEN_148 | _GEN_3826; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3836 = 2'h0 == opidx ? 32'h262b823 : _GEN_3827; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3837 = 2'h1 == opidx ? 32'h262b823 : _GEN_3828; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3838 = 2'h2 == opidx ? 32'h262b823 : _GEN_3829; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3839 = 2'h3 == opidx ? 32'h262b823 : _GEN_3830; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3840 = _GEN_1180 ? _cnt_T : _GEN_3831; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3841 = cnt[10] ? _GEN_3832 : _GEN_3823; // @[NulCtrlMP.scala 755:23]
  wire  _GEN_3842 = cnt[10] ? _GEN_3833 : _GEN_3824; // @[NulCtrlMP.scala 755:23]
  wire  _GEN_3843 = cnt[10] ? _GEN_3834 : _GEN_3825; // @[NulCtrlMP.scala 755:23]
  wire  _GEN_3844 = cnt[10] ? _GEN_3835 : _GEN_3826; // @[NulCtrlMP.scala 755:23]
  wire [31:0] _GEN_3845 = cnt[10] ? _GEN_3836 : _GEN_3827; // @[NulCtrlMP.scala 755:23]
  wire [31:0] _GEN_3846 = cnt[10] ? _GEN_3837 : _GEN_3828; // @[NulCtrlMP.scala 755:23]
  wire [31:0] _GEN_3847 = cnt[10] ? _GEN_3838 : _GEN_3829; // @[NulCtrlMP.scala 755:23]
  wire [31:0] _GEN_3848 = cnt[10] ? _GEN_3839 : _GEN_3830; // @[NulCtrlMP.scala 755:23]
  wire [128:0] _GEN_3849 = cnt[10] ? _GEN_3840 : _GEN_3831; // @[NulCtrlMP.scala 755:23]
  wire  _GEN_3850 = _GEN_145 | _GEN_3841; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3851 = _GEN_146 | _GEN_3842; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3852 = _GEN_147 | _GEN_3843; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3853 = _GEN_148 | _GEN_3844; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3854 = 2'h0 == opidx ? 32'h262bc23 : _GEN_3845; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3855 = 2'h1 == opidx ? 32'h262bc23 : _GEN_3846; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3856 = 2'h2 == opidx ? 32'h262bc23 : _GEN_3847; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3857 = 2'h3 == opidx ? 32'h262bc23 : _GEN_3848; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3858 = _GEN_1180 ? _cnt_T : _GEN_3849; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3859 = cnt[11] ? _GEN_3850 : _GEN_3841; // @[NulCtrlMP.scala 756:23]
  wire  _GEN_3860 = cnt[11] ? _GEN_3851 : _GEN_3842; // @[NulCtrlMP.scala 756:23]
  wire  _GEN_3861 = cnt[11] ? _GEN_3852 : _GEN_3843; // @[NulCtrlMP.scala 756:23]
  wire  _GEN_3862 = cnt[11] ? _GEN_3853 : _GEN_3844; // @[NulCtrlMP.scala 756:23]
  wire [31:0] _GEN_3863 = cnt[11] ? _GEN_3854 : _GEN_3845; // @[NulCtrlMP.scala 756:23]
  wire [31:0] _GEN_3864 = cnt[11] ? _GEN_3855 : _GEN_3846; // @[NulCtrlMP.scala 756:23]
  wire [31:0] _GEN_3865 = cnt[11] ? _GEN_3856 : _GEN_3847; // @[NulCtrlMP.scala 756:23]
  wire [31:0] _GEN_3866 = cnt[11] ? _GEN_3857 : _GEN_3848; // @[NulCtrlMP.scala 756:23]
  wire [128:0] _GEN_3867 = cnt[11] ? _GEN_3858 : _GEN_3849; // @[NulCtrlMP.scala 756:23]
  wire  _GEN_3868 = _GEN_145 | _GEN_3859; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3869 = _GEN_146 | _GEN_3860; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3870 = _GEN_147 | _GEN_3861; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3871 = _GEN_148 | _GEN_3862; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3872 = 2'h0 == opidx ? 32'h4028293 : _GEN_3863; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3873 = 2'h1 == opidx ? 32'h4028293 : _GEN_3864; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3874 = 2'h2 == opidx ? 32'h4028293 : _GEN_3865; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3875 = 2'h3 == opidx ? 32'h4028293 : _GEN_3866; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3876 = _GEN_1180 ? _cnt_T : _GEN_3867; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3877 = cnt[12] ? _GEN_3868 : _GEN_3859; // @[NulCtrlMP.scala 757:23]
  wire  _GEN_3878 = cnt[12] ? _GEN_3869 : _GEN_3860; // @[NulCtrlMP.scala 757:23]
  wire  _GEN_3879 = cnt[12] ? _GEN_3870 : _GEN_3861; // @[NulCtrlMP.scala 757:23]
  wire  _GEN_3880 = cnt[12] ? _GEN_3871 : _GEN_3862; // @[NulCtrlMP.scala 757:23]
  wire [31:0] _GEN_3881 = cnt[12] ? _GEN_3872 : _GEN_3863; // @[NulCtrlMP.scala 757:23]
  wire [31:0] _GEN_3882 = cnt[12] ? _GEN_3873 : _GEN_3864; // @[NulCtrlMP.scala 757:23]
  wire [31:0] _GEN_3883 = cnt[12] ? _GEN_3874 : _GEN_3865; // @[NulCtrlMP.scala 757:23]
  wire [31:0] _GEN_3884 = cnt[12] ? _GEN_3875 : _GEN_3866; // @[NulCtrlMP.scala 757:23]
  wire [128:0] _GEN_3885 = cnt[12] ? _GEN_3876 : _GEN_3867; // @[NulCtrlMP.scala 757:23]
  wire  _GEN_3886 = _GEN_145 | _GEN_3627; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3887 = _GEN_146 | _GEN_3628; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3888 = _GEN_147 | _GEN_3629; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3889 = _GEN_148 | _GEN_3630; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_3890 = ~_GEN_1252 ? _cnt_T : _GEN_3885; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_3891 = cnt[13] ? _GEN_3886 : _GEN_3627; // @[NulCtrlMP.scala 758:23]
  wire  _GEN_3892 = cnt[13] ? _GEN_3887 : _GEN_3628; // @[NulCtrlMP.scala 758:23]
  wire  _GEN_3893 = cnt[13] ? _GEN_3888 : _GEN_3629; // @[NulCtrlMP.scala 758:23]
  wire  _GEN_3894 = cnt[13] ? _GEN_3889 : _GEN_3630; // @[NulCtrlMP.scala 758:23]
  wire [128:0] _GEN_3895 = cnt[13] ? _GEN_3890 : _GEN_3885; // @[NulCtrlMP.scala 758:23]
  wire [7:0] _pg_loop_cnt_T_1 = pg_loop_cnt + 8'h1; // @[NulCtrlMP.scala 762:44]
  wire [128:0] _GEN_3896 = pg_loop_cnt != 8'h3f ? 129'h10 : _cnt_T; // @[NulCtrlMP.scala 760:40 761:21 764:21]
  wire [7:0] _GEN_3897 = pg_loop_cnt != 8'h3f ? _pg_loop_cnt_T_1 : 8'h0; // @[NulCtrlMP.scala 760:40 762:29 765:29]
  wire [128:0] _GEN_3898 = cnt[14] ? _GEN_3896 : _GEN_3895; // @[NulCtrlMP.scala 759:23]
  wire [7:0] _GEN_3899 = cnt[14] ? _GEN_3897 : pg_loop_cnt; // @[NulCtrlMP.scala 759:23 742:30]
  wire  _GEN_3900 = _GEN_145 | _GEN_3877; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3901 = _GEN_146 | _GEN_3878; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3902 = _GEN_147 | _GEN_3879; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_3903 = _GEN_148 | _GEN_3880; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_3904 = 2'h0 == opidx ? 32'h330000f : _GEN_3881; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3905 = 2'h1 == opidx ? 32'h330000f : _GEN_3882; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3906 = 2'h2 == opidx ? 32'h330000f : _GEN_3883; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_3907 = 2'h3 == opidx ? 32'h330000f : _GEN_3884; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_3908 = _GEN_1180 ? _cnt_T : _GEN_3898; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_3909 = cnt[15] ? _GEN_3900 : _GEN_3877; // @[NulCtrlMP.scala 768:23]
  wire  _GEN_3910 = cnt[15] ? _GEN_3901 : _GEN_3878; // @[NulCtrlMP.scala 768:23]
  wire  _GEN_3911 = cnt[15] ? _GEN_3902 : _GEN_3879; // @[NulCtrlMP.scala 768:23]
  wire  _GEN_3912 = cnt[15] ? _GEN_3903 : _GEN_3880; // @[NulCtrlMP.scala 768:23]
  wire [31:0] _GEN_3913 = cnt[15] ? _GEN_3904 : _GEN_3881; // @[NulCtrlMP.scala 768:23]
  wire [31:0] _GEN_3914 = cnt[15] ? _GEN_3905 : _GEN_3882; // @[NulCtrlMP.scala 768:23]
  wire [31:0] _GEN_3915 = cnt[15] ? _GEN_3906 : _GEN_3883; // @[NulCtrlMP.scala 768:23]
  wire [31:0] _GEN_3916 = cnt[15] ? _GEN_3907 : _GEN_3884; // @[NulCtrlMP.scala 768:23]
  wire [128:0] _GEN_3917 = cnt[15] ? _GEN_3908 : _GEN_3898; // @[NulCtrlMP.scala 768:23]
  wire  _GEN_3918 = _GEN_145 | _GEN_3891; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3919 = _GEN_146 | _GEN_3892; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3920 = _GEN_147 | _GEN_3893; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_3921 = _GEN_148 | _GEN_3894; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_3922 = ~_GEN_1252 ? _cnt_T : _GEN_3917; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_3923 = cnt[16] ? _GEN_3918 : _GEN_3891; // @[NulCtrlMP.scala 769:23]
  wire  _GEN_3924 = cnt[16] ? _GEN_3919 : _GEN_3892; // @[NulCtrlMP.scala 769:23]
  wire  _GEN_3925 = cnt[16] ? _GEN_3920 : _GEN_3893; // @[NulCtrlMP.scala 769:23]
  wire  _GEN_3926 = cnt[16] ? _GEN_3921 : _GEN_3894; // @[NulCtrlMP.scala 769:23]
  wire [128:0] _GEN_3927 = cnt[16] ? _GEN_3922 : _GEN_3917; // @[NulCtrlMP.scala 769:23]
  wire  _GEN_3928 = _GEN_145 | _GEN_3711; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3929 = _GEN_146 | _GEN_3712; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3930 = _GEN_147 | _GEN_3713; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3931 = _GEN_148 | _GEN_3714; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_3932 = 2'h0 == opidx ? 5'h5 : _GEN_3715; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3933 = 2'h1 == opidx ? 5'h5 : _GEN_3716; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3934 = 2'h2 == opidx ? 5'h5 : _GEN_3717; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3935 = 2'h3 == opidx ? 5'h5 : _GEN_3718; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_3936 = 2'h0 == opidx ? regback_0 : _GEN_3719; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3937 = 2'h1 == opidx ? regback_0 : _GEN_3720; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3938 = 2'h2 == opidx ? regback_0 : _GEN_3721; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3939 = 2'h3 == opidx ? regback_0 : _GEN_3722; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_3940 = ~_GEN_1128 ? _cnt_T : _GEN_3927; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_3941 = cnt[17] ? _GEN_3928 : _GEN_3711; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3942 = cnt[17] ? _GEN_3929 : _GEN_3712; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3943 = cnt[17] ? _GEN_3930 : _GEN_3713; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3944 = cnt[17] ? _GEN_3931 : _GEN_3714; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3945 = cnt[17] ? _GEN_3932 : _GEN_3715; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3946 = cnt[17] ? _GEN_3933 : _GEN_3716; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3947 = cnt[17] ? _GEN_3934 : _GEN_3717; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3948 = cnt[17] ? _GEN_3935 : _GEN_3718; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3949 = cnt[17] ? _GEN_3936 : _GEN_3719; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3950 = cnt[17] ? _GEN_3937 : _GEN_3720; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3951 = cnt[17] ? _GEN_3938 : _GEN_3721; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3952 = cnt[17] ? _GEN_3939 : _GEN_3722; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3953 = cnt[17] ? _GEN_3940 : _GEN_3927; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3954 = _GEN_145 | _GEN_3941; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3955 = _GEN_146 | _GEN_3942; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3956 = _GEN_147 | _GEN_3943; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_3957 = _GEN_148 | _GEN_3944; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_3958 = 2'h0 == opidx ? 5'h6 : _GEN_3945; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3959 = 2'h1 == opidx ? 5'h6 : _GEN_3946; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3960 = 2'h2 == opidx ? 5'h6 : _GEN_3947; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_3961 = 2'h3 == opidx ? 5'h6 : _GEN_3948; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_3962 = 2'h0 == opidx ? regback_1 : _GEN_3949; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3963 = 2'h1 == opidx ? regback_1 : _GEN_3950; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3964 = 2'h2 == opidx ? regback_1 : _GEN_3951; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_3965 = 2'h3 == opidx ? regback_1 : _GEN_3952; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_3966 = ~_GEN_1128 ? _cnt_T : _GEN_3953; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_3967 = cnt[18] ? _GEN_3954 : _GEN_3941; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3968 = cnt[18] ? _GEN_3955 : _GEN_3942; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3969 = cnt[18] ? _GEN_3956 : _GEN_3943; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_3970 = cnt[18] ? _GEN_3957 : _GEN_3944; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3971 = cnt[18] ? _GEN_3958 : _GEN_3945; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3972 = cnt[18] ? _GEN_3959 : _GEN_3946; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3973 = cnt[18] ? _GEN_3960 : _GEN_3947; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_3974 = cnt[18] ? _GEN_3961 : _GEN_3948; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3975 = cnt[18] ? _GEN_3962 : _GEN_3949; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3976 = cnt[18] ? _GEN_3963 : _GEN_3950; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3977 = cnt[18] ? _GEN_3964 : _GEN_3951; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_3978 = cnt[18] ? _GEN_3965 : _GEN_3952; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3979 = cnt[18] ? _GEN_3966 : _GEN_3953; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_3980 = cnt[19] ? 129'h1 : _GEN_3979; // @[NulCtrlMP.scala 771:23 772:17]
  wire [4:0] _GEN_3981 = cnt[19] ? 5'h5 : _GEN_3631; // @[NulCtrlMP.scala 771:23 773:19]
  wire  _GEN_3982 = state == 5'h13 ? _GEN_3662 : _GEN_3600; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_3983 = state == 5'h13 ? _GEN_3663 : _GEN_3601; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_3984 = state == 5'h13 ? _GEN_3664 : _GEN_3602; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_3985 = state == 5'h13 ? _GEN_3665 : _GEN_3603; // @[NulCtrlMP.scala 745:32]
  wire [4:0] _GEN_3986 = state == 5'h13 ? _GEN_3971 : _GEN_3604; // @[NulCtrlMP.scala 745:32]
  wire [4:0] _GEN_3987 = state == 5'h13 ? _GEN_3972 : _GEN_3605; // @[NulCtrlMP.scala 745:32]
  wire [4:0] _GEN_3988 = state == 5'h13 ? _GEN_3973 : _GEN_3606; // @[NulCtrlMP.scala 745:32]
  wire [4:0] _GEN_3989 = state == 5'h13 ? _GEN_3974 : _GEN_3607; // @[NulCtrlMP.scala 745:32]
  wire [128:0] _GEN_3990 = state == 5'h13 ? _GEN_3980 : _GEN_3608; // @[NulCtrlMP.scala 745:32]
  wire [63:0] _GEN_3991 = state == 5'h13 ? _GEN_3651 : _GEN_3609; // @[NulCtrlMP.scala 745:32]
  wire [63:0] _GEN_3992 = state == 5'h13 ? _GEN_3671 : _GEN_3610; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_3993 = state == 5'h13 ? _GEN_3967 : _GEN_3611; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_3994 = state == 5'h13 ? _GEN_3968 : _GEN_3612; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_3995 = state == 5'h13 ? _GEN_3969 : _GEN_3613; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_3996 = state == 5'h13 ? _GEN_3970 : _GEN_3614; // @[NulCtrlMP.scala 745:32]
  wire [63:0] _GEN_3997 = state == 5'h13 ? _GEN_3975 : _GEN_3615; // @[NulCtrlMP.scala 745:32]
  wire [63:0] _GEN_3998 = state == 5'h13 ? _GEN_3976 : _GEN_3616; // @[NulCtrlMP.scala 745:32]
  wire [63:0] _GEN_3999 = state == 5'h13 ? _GEN_3977 : _GEN_3617; // @[NulCtrlMP.scala 745:32]
  wire [63:0] _GEN_4000 = state == 5'h13 ? _GEN_3978 : _GEN_3618; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_4001 = state == 5'h13 ? _GEN_3909 : _GEN_3619; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_4002 = state == 5'h13 ? _GEN_3910 : _GEN_3620; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_4003 = state == 5'h13 ? _GEN_3911 : _GEN_3621; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_4004 = state == 5'h13 ? _GEN_3912 : _GEN_3622; // @[NulCtrlMP.scala 745:32]
  wire [31:0] _GEN_4005 = state == 5'h13 ? _GEN_3913 : _GEN_3623; // @[NulCtrlMP.scala 745:32]
  wire [31:0] _GEN_4006 = state == 5'h13 ? _GEN_3914 : _GEN_3624; // @[NulCtrlMP.scala 745:32]
  wire [31:0] _GEN_4007 = state == 5'h13 ? _GEN_3915 : _GEN_3625; // @[NulCtrlMP.scala 745:32]
  wire [31:0] _GEN_4008 = state == 5'h13 ? _GEN_3916 : _GEN_3626; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_4009 = state == 5'h13 ? _GEN_3923 : _GEN_3627; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_4010 = state == 5'h13 ? _GEN_3924 : _GEN_3628; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_4011 = state == 5'h13 ? _GEN_3925 : _GEN_3629; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_4012 = state == 5'h13 ? _GEN_3926 : _GEN_3630; // @[NulCtrlMP.scala 745:32]
  wire [7:0] _GEN_4013 = state == 5'h13 ? _GEN_3899 : pg_loop_cnt; // @[NulCtrlMP.scala 742:30 745:32]
  wire [4:0] _GEN_4014 = state == 5'h13 ? _GEN_3981 : _GEN_3631; // @[NulCtrlMP.scala 745:32]
  wire  _GEN_4015 = _GEN_145 | _GEN_3982; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4016 = _GEN_146 | _GEN_3983; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4017 = _GEN_147 | _GEN_3984; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4018 = _GEN_148 | _GEN_3985; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4019 = 2'h0 == opidx ? 5'h5 : _GEN_3986; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4020 = 2'h1 == opidx ? 5'h5 : _GEN_3987; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4021 = 2'h2 == opidx ? 5'h5 : _GEN_3988; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4022 = 2'h3 == opidx ? 5'h5 : _GEN_3989; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4023 = _T_122 ? _cnt_T : _GEN_3990; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4024 = _T_122 ? _GEN_1349 : _GEN_3991; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_4025 = cnt[0] ? _GEN_4015 : _GEN_3982; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4026 = cnt[0] ? _GEN_4016 : _GEN_3983; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4027 = cnt[0] ? _GEN_4017 : _GEN_3984; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4028 = cnt[0] ? _GEN_4018 : _GEN_3985; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4029 = cnt[0] ? _GEN_4019 : _GEN_3986; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4030 = cnt[0] ? _GEN_4020 : _GEN_3987; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4031 = cnt[0] ? _GEN_4021 : _GEN_3988; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4032 = cnt[0] ? _GEN_4022 : _GEN_3989; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4033 = cnt[0] ? _GEN_4023 : _GEN_3990; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4034 = cnt[0] ? _GEN_4024 : _GEN_3991; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4035 = _GEN_145 | _GEN_4025; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4036 = _GEN_146 | _GEN_4026; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4037 = _GEN_147 | _GEN_4027; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4038 = _GEN_148 | _GEN_4028; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4039 = 2'h0 == opidx ? 5'h6 : _GEN_4029; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4040 = 2'h1 == opidx ? 5'h6 : _GEN_4030; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4041 = 2'h2 == opidx ? 5'h6 : _GEN_4031; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4042 = 2'h3 == opidx ? 5'h6 : _GEN_4032; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4043 = _T_122 ? _cnt_T : _GEN_4033; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4044 = _T_122 ? _GEN_1349 : _GEN_3992; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_4045 = cnt[1] ? _GEN_4035 : _GEN_4025; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4046 = cnt[1] ? _GEN_4036 : _GEN_4026; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4047 = cnt[1] ? _GEN_4037 : _GEN_4027; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4048 = cnt[1] ? _GEN_4038 : _GEN_4028; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4049 = cnt[1] ? _GEN_4039 : _GEN_4029; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4050 = cnt[1] ? _GEN_4040 : _GEN_4030; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4051 = cnt[1] ? _GEN_4041 : _GEN_4031; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4052 = cnt[1] ? _GEN_4042 : _GEN_4032; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4053 = cnt[1] ? _GEN_4043 : _GEN_4033; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4054 = cnt[1] ? _GEN_4044 : _GEN_3992; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4055 = _GEN_145 | _GEN_4045; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4056 = _GEN_146 | _GEN_4046; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4057 = _GEN_147 | _GEN_4047; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4058 = _GEN_148 | _GEN_4048; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4059 = 2'h0 == opidx ? 5'h7 : _GEN_4049; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4060 = 2'h1 == opidx ? 5'h7 : _GEN_4050; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4061 = 2'h2 == opidx ? 5'h7 : _GEN_4051; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4062 = 2'h3 == opidx ? 5'h7 : _GEN_4052; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4063 = _T_122 ? _cnt_T : _GEN_4053; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4064 = _T_122 ? _GEN_1349 : _GEN_2439; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_4065 = cnt[2] ? _GEN_4055 : _GEN_4045; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4066 = cnt[2] ? _GEN_4056 : _GEN_4046; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4067 = cnt[2] ? _GEN_4057 : _GEN_4047; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4068 = cnt[2] ? _GEN_4058 : _GEN_4048; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4069 = cnt[2] ? _GEN_4059 : _GEN_4049; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4070 = cnt[2] ? _GEN_4060 : _GEN_4050; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4071 = cnt[2] ? _GEN_4061 : _GEN_4051; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4072 = cnt[2] ? _GEN_4062 : _GEN_4052; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4073 = cnt[2] ? _GEN_4063 : _GEN_4053; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4074 = cnt[2] ? _GEN_4064 : _GEN_2439; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4075 = _GEN_145 | _GEN_4065; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4076 = _GEN_146 | _GEN_4066; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4077 = _GEN_147 | _GEN_4067; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4078 = _GEN_148 | _GEN_4068; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4079 = 2'h0 == opidx ? 5'h8 : _GEN_4069; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4080 = 2'h1 == opidx ? 5'h8 : _GEN_4070; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4081 = 2'h2 == opidx ? 5'h8 : _GEN_4071; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4082 = 2'h3 == opidx ? 5'h8 : _GEN_4072; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4083 = _T_122 ? _cnt_T : _GEN_4073; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4084 = _T_122 ? _GEN_1349 : regback_3; // @[NulCtrlMP.scala 353:36 355:17 346:26]
  wire  _GEN_4085 = cnt[3] ? _GEN_4075 : _GEN_4065; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4086 = cnt[3] ? _GEN_4076 : _GEN_4066; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4087 = cnt[3] ? _GEN_4077 : _GEN_4067; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4088 = cnt[3] ? _GEN_4078 : _GEN_4068; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4089 = cnt[3] ? _GEN_4079 : _GEN_4069; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4090 = cnt[3] ? _GEN_4080 : _GEN_4070; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4091 = cnt[3] ? _GEN_4081 : _GEN_4071; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4092 = cnt[3] ? _GEN_4082 : _GEN_4072; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4093 = cnt[3] ? _GEN_4083 : _GEN_4073; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4094 = cnt[3] ? _GEN_4084 : regback_3; // @[NulCtrlMP.scala 346:26 408:32]
  wire  _GEN_4095 = _GEN_145 | _GEN_4085; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4096 = _GEN_146 | _GEN_4086; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4097 = _GEN_147 | _GEN_4087; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4098 = _GEN_148 | _GEN_4088; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4099 = 2'h0 == opidx ? 5'h9 : _GEN_4089; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4100 = 2'h1 == opidx ? 5'h9 : _GEN_4090; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4101 = 2'h2 == opidx ? 5'h9 : _GEN_4091; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4102 = 2'h3 == opidx ? 5'h9 : _GEN_4092; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4103 = _T_122 ? _cnt_T : _GEN_4093; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4104 = _T_122 ? _GEN_1349 : regback_4; // @[NulCtrlMP.scala 353:36 355:17 346:26]
  wire  _GEN_4105 = cnt[4] ? _GEN_4095 : _GEN_4085; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4106 = cnt[4] ? _GEN_4096 : _GEN_4086; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4107 = cnt[4] ? _GEN_4097 : _GEN_4087; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4108 = cnt[4] ? _GEN_4098 : _GEN_4088; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4109 = cnt[4] ? _GEN_4099 : _GEN_4089; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4110 = cnt[4] ? _GEN_4100 : _GEN_4090; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4111 = cnt[4] ? _GEN_4101 : _GEN_4091; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4112 = cnt[4] ? _GEN_4102 : _GEN_4092; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4113 = cnt[4] ? _GEN_4103 : _GEN_4093; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4114 = cnt[4] ? _GEN_4104 : regback_4; // @[NulCtrlMP.scala 346:26 408:32]
  wire  _GEN_4115 = _GEN_145 | _GEN_4105; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4116 = _GEN_146 | _GEN_4106; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4117 = _GEN_147 | _GEN_4107; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4118 = _GEN_148 | _GEN_4108; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4119 = 2'h0 == opidx ? 5'ha : _GEN_4109; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4120 = 2'h1 == opidx ? 5'ha : _GEN_4110; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4121 = 2'h2 == opidx ? 5'ha : _GEN_4111; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4122 = 2'h3 == opidx ? 5'ha : _GEN_4112; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4123 = _T_122 ? _cnt_T : _GEN_4113; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4124 = _T_122 ? _GEN_1349 : regback_5; // @[NulCtrlMP.scala 353:36 355:17 346:26]
  wire  _GEN_4125 = cnt[5] ? _GEN_4115 : _GEN_4105; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4126 = cnt[5] ? _GEN_4116 : _GEN_4106; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4127 = cnt[5] ? _GEN_4117 : _GEN_4107; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4128 = cnt[5] ? _GEN_4118 : _GEN_4108; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4129 = cnt[5] ? _GEN_4119 : _GEN_4109; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4130 = cnt[5] ? _GEN_4120 : _GEN_4110; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4131 = cnt[5] ? _GEN_4121 : _GEN_4111; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4132 = cnt[5] ? _GEN_4122 : _GEN_4112; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4133 = cnt[5] ? _GEN_4123 : _GEN_4113; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4134 = cnt[5] ? _GEN_4124 : regback_5; // @[NulCtrlMP.scala 346:26 408:32]
  wire  _GEN_4135 = _GEN_145 | _GEN_4125; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4136 = _GEN_146 | _GEN_4126; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4137 = _GEN_147 | _GEN_4127; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4138 = _GEN_148 | _GEN_4128; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4139 = 2'h0 == opidx ? 5'hb : _GEN_4129; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4140 = 2'h1 == opidx ? 5'hb : _GEN_4130; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4141 = 2'h2 == opidx ? 5'hb : _GEN_4131; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4142 = 2'h3 == opidx ? 5'hb : _GEN_4132; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4143 = _T_122 ? _cnt_T : _GEN_4133; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4144 = _T_122 ? _GEN_1349 : regback_6; // @[NulCtrlMP.scala 353:36 355:17 346:26]
  wire  _GEN_4145 = cnt[6] ? _GEN_4135 : _GEN_4125; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4146 = cnt[6] ? _GEN_4136 : _GEN_4126; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4147 = cnt[6] ? _GEN_4137 : _GEN_4127; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4148 = cnt[6] ? _GEN_4138 : _GEN_4128; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4149 = cnt[6] ? _GEN_4139 : _GEN_4129; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4150 = cnt[6] ? _GEN_4140 : _GEN_4130; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4151 = cnt[6] ? _GEN_4141 : _GEN_4131; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4152 = cnt[6] ? _GEN_4142 : _GEN_4132; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4153 = cnt[6] ? _GEN_4143 : _GEN_4133; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4154 = cnt[6] ? _GEN_4144 : regback_6; // @[NulCtrlMP.scala 346:26 408:32]
  wire  _GEN_4155 = _GEN_145 | _GEN_4145; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4156 = _GEN_146 | _GEN_4146; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4157 = _GEN_147 | _GEN_4147; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4158 = _GEN_148 | _GEN_4148; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4159 = 2'h0 == opidx ? 5'hc : _GEN_4149; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4160 = 2'h1 == opidx ? 5'hc : _GEN_4150; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4161 = 2'h2 == opidx ? 5'hc : _GEN_4151; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4162 = 2'h3 == opidx ? 5'hc : _GEN_4152; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4163 = _T_122 ? _cnt_T : _GEN_4153; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4164 = _T_122 ? _GEN_1349 : regback_7; // @[NulCtrlMP.scala 353:36 355:17 346:26]
  wire  _GEN_4165 = cnt[7] ? _GEN_4155 : _GEN_4145; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4166 = cnt[7] ? _GEN_4156 : _GEN_4146; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4167 = cnt[7] ? _GEN_4157 : _GEN_4147; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4168 = cnt[7] ? _GEN_4158 : _GEN_4148; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4169 = cnt[7] ? _GEN_4159 : _GEN_4149; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4170 = cnt[7] ? _GEN_4160 : _GEN_4150; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4171 = cnt[7] ? _GEN_4161 : _GEN_4151; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4172 = cnt[7] ? _GEN_4162 : _GEN_4152; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4173 = cnt[7] ? _GEN_4163 : _GEN_4153; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4174 = cnt[7] ? _GEN_4164 : regback_7; // @[NulCtrlMP.scala 346:26 408:32]
  wire  _GEN_4175 = _GEN_145 | _GEN_4165; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4176 = _GEN_146 | _GEN_4166; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4177 = _GEN_147 | _GEN_4167; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4178 = _GEN_148 | _GEN_4168; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4179 = 2'h0 == opidx ? 5'hd : _GEN_4169; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4180 = 2'h1 == opidx ? 5'hd : _GEN_4170; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4181 = 2'h2 == opidx ? 5'hd : _GEN_4171; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4182 = 2'h3 == opidx ? 5'hd : _GEN_4172; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4183 = _T_122 ? _cnt_T : _GEN_4173; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4184 = _T_122 ? _GEN_1349 : regback_8; // @[NulCtrlMP.scala 353:36 355:17 346:26]
  wire  _GEN_4185 = cnt[8] ? _GEN_4175 : _GEN_4165; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4186 = cnt[8] ? _GEN_4176 : _GEN_4166; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4187 = cnt[8] ? _GEN_4177 : _GEN_4167; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4188 = cnt[8] ? _GEN_4178 : _GEN_4168; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4189 = cnt[8] ? _GEN_4179 : _GEN_4169; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4190 = cnt[8] ? _GEN_4180 : _GEN_4170; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4191 = cnt[8] ? _GEN_4181 : _GEN_4171; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4192 = cnt[8] ? _GEN_4182 : _GEN_4172; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4193 = cnt[8] ? _GEN_4183 : _GEN_4173; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4194 = cnt[8] ? _GEN_4184 : regback_8; // @[NulCtrlMP.scala 346:26 408:32]
  wire  _GEN_4195 = _GEN_145 | _GEN_4185; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4196 = _GEN_146 | _GEN_4186; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4197 = _GEN_147 | _GEN_4187; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4198 = _GEN_148 | _GEN_4188; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4199 = 2'h0 == opidx ? 5'he : _GEN_4189; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4200 = 2'h1 == opidx ? 5'he : _GEN_4190; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4201 = 2'h2 == opidx ? 5'he : _GEN_4191; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4202 = 2'h3 == opidx ? 5'he : _GEN_4192; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4203 = _T_122 ? _cnt_T : _GEN_4193; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_4205 = cnt[9] ? _GEN_4195 : _GEN_4185; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4206 = cnt[9] ? _GEN_4196 : _GEN_4186; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4207 = cnt[9] ? _GEN_4197 : _GEN_4187; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4208 = cnt[9] ? _GEN_4198 : _GEN_4188; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4209 = cnt[9] ? _GEN_4199 : _GEN_4189; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4210 = cnt[9] ? _GEN_4200 : _GEN_4190; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4211 = cnt[9] ? _GEN_4201 : _GEN_4191; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4212 = cnt[9] ? _GEN_4202 : _GEN_4192; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4213 = cnt[9] ? _GEN_4203 : _GEN_4193; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4215 = _GEN_145 | _GEN_3993; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4216 = _GEN_146 | _GEN_3994; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4217 = _GEN_147 | _GEN_3995; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4218 = _GEN_148 | _GEN_3996; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4219 = 2'h0 == opidx ? 5'h5 : _GEN_4209; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4220 = 2'h1 == opidx ? 5'h5 : _GEN_4210; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4221 = 2'h2 == opidx ? 5'h5 : _GEN_4211; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4222 = 2'h3 == opidx ? 5'h5 : _GEN_4212; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4223 = 2'h0 == opidx ? pg_base_addr7 : _GEN_3997; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4224 = 2'h1 == opidx ? pg_base_addr7 : _GEN_3998; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4225 = 2'h2 == opidx ? pg_base_addr7 : _GEN_3999; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4226 = 2'h3 == opidx ? pg_base_addr7 : _GEN_4000; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4227 = ~_GEN_1128 ? _cnt_T : _GEN_4213; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4228 = cnt[10] ? _GEN_4215 : _GEN_3993; // @[NulCtrlMP.scala 779:23]
  wire  _GEN_4229 = cnt[10] ? _GEN_4216 : _GEN_3994; // @[NulCtrlMP.scala 779:23]
  wire  _GEN_4230 = cnt[10] ? _GEN_4217 : _GEN_3995; // @[NulCtrlMP.scala 779:23]
  wire  _GEN_4231 = cnt[10] ? _GEN_4218 : _GEN_3996; // @[NulCtrlMP.scala 779:23]
  wire [4:0] _GEN_4232 = cnt[10] ? _GEN_4219 : _GEN_4209; // @[NulCtrlMP.scala 779:23]
  wire [4:0] _GEN_4233 = cnt[10] ? _GEN_4220 : _GEN_4210; // @[NulCtrlMP.scala 779:23]
  wire [4:0] _GEN_4234 = cnt[10] ? _GEN_4221 : _GEN_4211; // @[NulCtrlMP.scala 779:23]
  wire [4:0] _GEN_4235 = cnt[10] ? _GEN_4222 : _GEN_4212; // @[NulCtrlMP.scala 779:23]
  wire [63:0] _GEN_4236 = cnt[10] ? _GEN_4223 : _GEN_3997; // @[NulCtrlMP.scala 779:23]
  wire [63:0] _GEN_4237 = cnt[10] ? _GEN_4224 : _GEN_3998; // @[NulCtrlMP.scala 779:23]
  wire [63:0] _GEN_4238 = cnt[10] ? _GEN_4225 : _GEN_3999; // @[NulCtrlMP.scala 779:23]
  wire [63:0] _GEN_4239 = cnt[10] ? _GEN_4226 : _GEN_4000; // @[NulCtrlMP.scala 779:23]
  wire [128:0] _GEN_4240 = cnt[10] ? _GEN_4227 : _GEN_4213; // @[NulCtrlMP.scala 779:23]
  wire  _GEN_4241 = _GEN_145 | _GEN_4228; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4242 = _GEN_146 | _GEN_4229; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4243 = _GEN_147 | _GEN_4230; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4244 = _GEN_148 | _GEN_4231; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4245 = 2'h0 == opidx ? 5'he : _GEN_4232; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4246 = 2'h1 == opidx ? 5'he : _GEN_4233; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4247 = 2'h2 == opidx ? 5'he : _GEN_4234; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4248 = 2'h3 == opidx ? 5'he : _GEN_4235; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4249 = 2'h0 == opidx ? pg_base_addr2 : _GEN_4236; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4250 = 2'h1 == opidx ? pg_base_addr2 : _GEN_4237; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4251 = 2'h2 == opidx ? pg_base_addr2 : _GEN_4238; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4252 = 2'h3 == opidx ? pg_base_addr2 : _GEN_4239; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4253 = ~_GEN_1128 ? _cnt_T : _GEN_4240; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4254 = cnt[11] ? _GEN_4241 : _GEN_4228; // @[NulCtrlMP.scala 780:23]
  wire  _GEN_4255 = cnt[11] ? _GEN_4242 : _GEN_4229; // @[NulCtrlMP.scala 780:23]
  wire  _GEN_4256 = cnt[11] ? _GEN_4243 : _GEN_4230; // @[NulCtrlMP.scala 780:23]
  wire  _GEN_4257 = cnt[11] ? _GEN_4244 : _GEN_4231; // @[NulCtrlMP.scala 780:23]
  wire [4:0] _GEN_4258 = cnt[11] ? _GEN_4245 : _GEN_4232; // @[NulCtrlMP.scala 780:23]
  wire [4:0] _GEN_4259 = cnt[11] ? _GEN_4246 : _GEN_4233; // @[NulCtrlMP.scala 780:23]
  wire [4:0] _GEN_4260 = cnt[11] ? _GEN_4247 : _GEN_4234; // @[NulCtrlMP.scala 780:23]
  wire [4:0] _GEN_4261 = cnt[11] ? _GEN_4248 : _GEN_4235; // @[NulCtrlMP.scala 780:23]
  wire [63:0] _GEN_4262 = cnt[11] ? _GEN_4249 : _GEN_4236; // @[NulCtrlMP.scala 780:23]
  wire [63:0] _GEN_4263 = cnt[11] ? _GEN_4250 : _GEN_4237; // @[NulCtrlMP.scala 780:23]
  wire [63:0] _GEN_4264 = cnt[11] ? _GEN_4251 : _GEN_4238; // @[NulCtrlMP.scala 780:23]
  wire [63:0] _GEN_4265 = cnt[11] ? _GEN_4252 : _GEN_4239; // @[NulCtrlMP.scala 780:23]
  wire [128:0] _GEN_4266 = cnt[11] ? _GEN_4253 : _GEN_4240; // @[NulCtrlMP.scala 780:23]
  wire  _GEN_4267 = _GEN_145 | _GEN_4001; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4268 = _GEN_146 | _GEN_4002; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4269 = _GEN_147 | _GEN_4003; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4270 = _GEN_148 | _GEN_4004; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4271 = 2'h0 == opidx ? 32'h2b303 : _GEN_4005; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4272 = 2'h1 == opidx ? 32'h2b303 : _GEN_4006; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4273 = 2'h2 == opidx ? 32'h2b303 : _GEN_4007; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4274 = 2'h3 == opidx ? 32'h2b303 : _GEN_4008; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4275 = _GEN_1180 ? _cnt_T : _GEN_4266; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4276 = cnt[12] ? _GEN_4267 : _GEN_4001; // @[NulCtrlMP.scala 781:23]
  wire  _GEN_4277 = cnt[12] ? _GEN_4268 : _GEN_4002; // @[NulCtrlMP.scala 781:23]
  wire  _GEN_4278 = cnt[12] ? _GEN_4269 : _GEN_4003; // @[NulCtrlMP.scala 781:23]
  wire  _GEN_4279 = cnt[12] ? _GEN_4270 : _GEN_4004; // @[NulCtrlMP.scala 781:23]
  wire [31:0] _GEN_4280 = cnt[12] ? _GEN_4271 : _GEN_4005; // @[NulCtrlMP.scala 781:23]
  wire [31:0] _GEN_4281 = cnt[12] ? _GEN_4272 : _GEN_4006; // @[NulCtrlMP.scala 781:23]
  wire [31:0] _GEN_4282 = cnt[12] ? _GEN_4273 : _GEN_4007; // @[NulCtrlMP.scala 781:23]
  wire [31:0] _GEN_4283 = cnt[12] ? _GEN_4274 : _GEN_4008; // @[NulCtrlMP.scala 781:23]
  wire [128:0] _GEN_4284 = cnt[12] ? _GEN_4275 : _GEN_4266; // @[NulCtrlMP.scala 781:23]
  wire  _GEN_4285 = _GEN_145 | _GEN_4276; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4286 = _GEN_146 | _GEN_4277; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4287 = _GEN_147 | _GEN_4278; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4288 = _GEN_148 | _GEN_4279; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4289 = 2'h0 == opidx ? 32'h82b383 : _GEN_4280; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4290 = 2'h1 == opidx ? 32'h82b383 : _GEN_4281; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4291 = 2'h2 == opidx ? 32'h82b383 : _GEN_4282; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4292 = 2'h3 == opidx ? 32'h82b383 : _GEN_4283; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4293 = _GEN_1180 ? _cnt_T : _GEN_4284; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4294 = cnt[13] ? _GEN_4285 : _GEN_4276; // @[NulCtrlMP.scala 782:23]
  wire  _GEN_4295 = cnt[13] ? _GEN_4286 : _GEN_4277; // @[NulCtrlMP.scala 782:23]
  wire  _GEN_4296 = cnt[13] ? _GEN_4287 : _GEN_4278; // @[NulCtrlMP.scala 782:23]
  wire  _GEN_4297 = cnt[13] ? _GEN_4288 : _GEN_4279; // @[NulCtrlMP.scala 782:23]
  wire [31:0] _GEN_4298 = cnt[13] ? _GEN_4289 : _GEN_4280; // @[NulCtrlMP.scala 782:23]
  wire [31:0] _GEN_4299 = cnt[13] ? _GEN_4290 : _GEN_4281; // @[NulCtrlMP.scala 782:23]
  wire [31:0] _GEN_4300 = cnt[13] ? _GEN_4291 : _GEN_4282; // @[NulCtrlMP.scala 782:23]
  wire [31:0] _GEN_4301 = cnt[13] ? _GEN_4292 : _GEN_4283; // @[NulCtrlMP.scala 782:23]
  wire [128:0] _GEN_4302 = cnt[13] ? _GEN_4293 : _GEN_4284; // @[NulCtrlMP.scala 782:23]
  wire  _GEN_4303 = _GEN_145 | _GEN_4294; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4304 = _GEN_146 | _GEN_4295; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4305 = _GEN_147 | _GEN_4296; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4306 = _GEN_148 | _GEN_4297; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4307 = 2'h0 == opidx ? 32'h102b403 : _GEN_4298; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4308 = 2'h1 == opidx ? 32'h102b403 : _GEN_4299; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4309 = 2'h2 == opidx ? 32'h102b403 : _GEN_4300; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4310 = 2'h3 == opidx ? 32'h102b403 : _GEN_4301; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4311 = _GEN_1180 ? _cnt_T : _GEN_4302; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4312 = cnt[14] ? _GEN_4303 : _GEN_4294; // @[NulCtrlMP.scala 783:23]
  wire  _GEN_4313 = cnt[14] ? _GEN_4304 : _GEN_4295; // @[NulCtrlMP.scala 783:23]
  wire  _GEN_4314 = cnt[14] ? _GEN_4305 : _GEN_4296; // @[NulCtrlMP.scala 783:23]
  wire  _GEN_4315 = cnt[14] ? _GEN_4306 : _GEN_4297; // @[NulCtrlMP.scala 783:23]
  wire [31:0] _GEN_4316 = cnt[14] ? _GEN_4307 : _GEN_4298; // @[NulCtrlMP.scala 783:23]
  wire [31:0] _GEN_4317 = cnt[14] ? _GEN_4308 : _GEN_4299; // @[NulCtrlMP.scala 783:23]
  wire [31:0] _GEN_4318 = cnt[14] ? _GEN_4309 : _GEN_4300; // @[NulCtrlMP.scala 783:23]
  wire [31:0] _GEN_4319 = cnt[14] ? _GEN_4310 : _GEN_4301; // @[NulCtrlMP.scala 783:23]
  wire [128:0] _GEN_4320 = cnt[14] ? _GEN_4311 : _GEN_4302; // @[NulCtrlMP.scala 783:23]
  wire  _GEN_4321 = _GEN_145 | _GEN_4312; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4322 = _GEN_146 | _GEN_4313; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4323 = _GEN_147 | _GEN_4314; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4324 = _GEN_148 | _GEN_4315; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4325 = 2'h0 == opidx ? 32'h182b483 : _GEN_4316; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4326 = 2'h1 == opidx ? 32'h182b483 : _GEN_4317; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4327 = 2'h2 == opidx ? 32'h182b483 : _GEN_4318; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4328 = 2'h3 == opidx ? 32'h182b483 : _GEN_4319; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4329 = _GEN_1180 ? _cnt_T : _GEN_4320; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4330 = cnt[15] ? _GEN_4321 : _GEN_4312; // @[NulCtrlMP.scala 784:23]
  wire  _GEN_4331 = cnt[15] ? _GEN_4322 : _GEN_4313; // @[NulCtrlMP.scala 784:23]
  wire  _GEN_4332 = cnt[15] ? _GEN_4323 : _GEN_4314; // @[NulCtrlMP.scala 784:23]
  wire  _GEN_4333 = cnt[15] ? _GEN_4324 : _GEN_4315; // @[NulCtrlMP.scala 784:23]
  wire [31:0] _GEN_4334 = cnt[15] ? _GEN_4325 : _GEN_4316; // @[NulCtrlMP.scala 784:23]
  wire [31:0] _GEN_4335 = cnt[15] ? _GEN_4326 : _GEN_4317; // @[NulCtrlMP.scala 784:23]
  wire [31:0] _GEN_4336 = cnt[15] ? _GEN_4327 : _GEN_4318; // @[NulCtrlMP.scala 784:23]
  wire [31:0] _GEN_4337 = cnt[15] ? _GEN_4328 : _GEN_4319; // @[NulCtrlMP.scala 784:23]
  wire [128:0] _GEN_4338 = cnt[15] ? _GEN_4329 : _GEN_4320; // @[NulCtrlMP.scala 784:23]
  wire  _GEN_4339 = _GEN_145 | _GEN_4330; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4340 = _GEN_146 | _GEN_4331; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4341 = _GEN_147 | _GEN_4332; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4342 = _GEN_148 | _GEN_4333; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4343 = 2'h0 == opidx ? 32'h202b503 : _GEN_4334; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4344 = 2'h1 == opidx ? 32'h202b503 : _GEN_4335; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4345 = 2'h2 == opidx ? 32'h202b503 : _GEN_4336; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4346 = 2'h3 == opidx ? 32'h202b503 : _GEN_4337; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4347 = _GEN_1180 ? _cnt_T : _GEN_4338; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4348 = cnt[16] ? _GEN_4339 : _GEN_4330; // @[NulCtrlMP.scala 785:23]
  wire  _GEN_4349 = cnt[16] ? _GEN_4340 : _GEN_4331; // @[NulCtrlMP.scala 785:23]
  wire  _GEN_4350 = cnt[16] ? _GEN_4341 : _GEN_4332; // @[NulCtrlMP.scala 785:23]
  wire  _GEN_4351 = cnt[16] ? _GEN_4342 : _GEN_4333; // @[NulCtrlMP.scala 785:23]
  wire [31:0] _GEN_4352 = cnt[16] ? _GEN_4343 : _GEN_4334; // @[NulCtrlMP.scala 785:23]
  wire [31:0] _GEN_4353 = cnt[16] ? _GEN_4344 : _GEN_4335; // @[NulCtrlMP.scala 785:23]
  wire [31:0] _GEN_4354 = cnt[16] ? _GEN_4345 : _GEN_4336; // @[NulCtrlMP.scala 785:23]
  wire [31:0] _GEN_4355 = cnt[16] ? _GEN_4346 : _GEN_4337; // @[NulCtrlMP.scala 785:23]
  wire [128:0] _GEN_4356 = cnt[16] ? _GEN_4347 : _GEN_4338; // @[NulCtrlMP.scala 785:23]
  wire  _GEN_4357 = _GEN_145 | _GEN_4348; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4358 = _GEN_146 | _GEN_4349; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4359 = _GEN_147 | _GEN_4350; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4360 = _GEN_148 | _GEN_4351; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4361 = 2'h0 == opidx ? 32'h282b583 : _GEN_4352; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4362 = 2'h1 == opidx ? 32'h282b583 : _GEN_4353; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4363 = 2'h2 == opidx ? 32'h282b583 : _GEN_4354; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4364 = 2'h3 == opidx ? 32'h282b583 : _GEN_4355; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4365 = _GEN_1180 ? _cnt_T : _GEN_4356; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4366 = cnt[17] ? _GEN_4357 : _GEN_4348; // @[NulCtrlMP.scala 786:23]
  wire  _GEN_4367 = cnt[17] ? _GEN_4358 : _GEN_4349; // @[NulCtrlMP.scala 786:23]
  wire  _GEN_4368 = cnt[17] ? _GEN_4359 : _GEN_4350; // @[NulCtrlMP.scala 786:23]
  wire  _GEN_4369 = cnt[17] ? _GEN_4360 : _GEN_4351; // @[NulCtrlMP.scala 786:23]
  wire [31:0] _GEN_4370 = cnt[17] ? _GEN_4361 : _GEN_4352; // @[NulCtrlMP.scala 786:23]
  wire [31:0] _GEN_4371 = cnt[17] ? _GEN_4362 : _GEN_4353; // @[NulCtrlMP.scala 786:23]
  wire [31:0] _GEN_4372 = cnt[17] ? _GEN_4363 : _GEN_4354; // @[NulCtrlMP.scala 786:23]
  wire [31:0] _GEN_4373 = cnt[17] ? _GEN_4364 : _GEN_4355; // @[NulCtrlMP.scala 786:23]
  wire [128:0] _GEN_4374 = cnt[17] ? _GEN_4365 : _GEN_4356; // @[NulCtrlMP.scala 786:23]
  wire  _GEN_4375 = _GEN_145 | _GEN_4366; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4376 = _GEN_146 | _GEN_4367; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4377 = _GEN_147 | _GEN_4368; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4378 = _GEN_148 | _GEN_4369; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4379 = 2'h0 == opidx ? 32'h302b603 : _GEN_4370; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4380 = 2'h1 == opidx ? 32'h302b603 : _GEN_4371; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4381 = 2'h2 == opidx ? 32'h302b603 : _GEN_4372; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4382 = 2'h3 == opidx ? 32'h302b603 : _GEN_4373; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4383 = _GEN_1180 ? _cnt_T : _GEN_4374; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4384 = cnt[18] ? _GEN_4375 : _GEN_4366; // @[NulCtrlMP.scala 787:23]
  wire  _GEN_4385 = cnt[18] ? _GEN_4376 : _GEN_4367; // @[NulCtrlMP.scala 787:23]
  wire  _GEN_4386 = cnt[18] ? _GEN_4377 : _GEN_4368; // @[NulCtrlMP.scala 787:23]
  wire  _GEN_4387 = cnt[18] ? _GEN_4378 : _GEN_4369; // @[NulCtrlMP.scala 787:23]
  wire [31:0] _GEN_4388 = cnt[18] ? _GEN_4379 : _GEN_4370; // @[NulCtrlMP.scala 787:23]
  wire [31:0] _GEN_4389 = cnt[18] ? _GEN_4380 : _GEN_4371; // @[NulCtrlMP.scala 787:23]
  wire [31:0] _GEN_4390 = cnt[18] ? _GEN_4381 : _GEN_4372; // @[NulCtrlMP.scala 787:23]
  wire [31:0] _GEN_4391 = cnt[18] ? _GEN_4382 : _GEN_4373; // @[NulCtrlMP.scala 787:23]
  wire [128:0] _GEN_4392 = cnt[18] ? _GEN_4383 : _GEN_4374; // @[NulCtrlMP.scala 787:23]
  wire  _GEN_4393 = _GEN_145 | _GEN_4384; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4394 = _GEN_146 | _GEN_4385; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4395 = _GEN_147 | _GEN_4386; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4396 = _GEN_148 | _GEN_4387; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4397 = 2'h0 == opidx ? 32'h382b683 : _GEN_4388; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4398 = 2'h1 == opidx ? 32'h382b683 : _GEN_4389; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4399 = 2'h2 == opidx ? 32'h382b683 : _GEN_4390; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4400 = 2'h3 == opidx ? 32'h382b683 : _GEN_4391; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4401 = _GEN_1180 ? _cnt_T : _GEN_4392; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4402 = cnt[19] ? _GEN_4393 : _GEN_4384; // @[NulCtrlMP.scala 788:23]
  wire  _GEN_4403 = cnt[19] ? _GEN_4394 : _GEN_4385; // @[NulCtrlMP.scala 788:23]
  wire  _GEN_4404 = cnt[19] ? _GEN_4395 : _GEN_4386; // @[NulCtrlMP.scala 788:23]
  wire  _GEN_4405 = cnt[19] ? _GEN_4396 : _GEN_4387; // @[NulCtrlMP.scala 788:23]
  wire [31:0] _GEN_4406 = cnt[19] ? _GEN_4397 : _GEN_4388; // @[NulCtrlMP.scala 788:23]
  wire [31:0] _GEN_4407 = cnt[19] ? _GEN_4398 : _GEN_4389; // @[NulCtrlMP.scala 788:23]
  wire [31:0] _GEN_4408 = cnt[19] ? _GEN_4399 : _GEN_4390; // @[NulCtrlMP.scala 788:23]
  wire [31:0] _GEN_4409 = cnt[19] ? _GEN_4400 : _GEN_4391; // @[NulCtrlMP.scala 788:23]
  wire [128:0] _GEN_4410 = cnt[19] ? _GEN_4401 : _GEN_4392; // @[NulCtrlMP.scala 788:23]
  wire  _GEN_4411 = _GEN_145 | _GEN_4402; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4412 = _GEN_146 | _GEN_4403; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4413 = _GEN_147 | _GEN_4404; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4414 = _GEN_148 | _GEN_4405; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4415 = 2'h0 == opidx ? 32'h673023 : _GEN_4406; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4416 = 2'h1 == opidx ? 32'h673023 : _GEN_4407; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4417 = 2'h2 == opidx ? 32'h673023 : _GEN_4408; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4418 = 2'h3 == opidx ? 32'h673023 : _GEN_4409; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4419 = _GEN_1180 ? _cnt_T : _GEN_4410; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4420 = cnt[20] ? _GEN_4411 : _GEN_4402; // @[NulCtrlMP.scala 789:23]
  wire  _GEN_4421 = cnt[20] ? _GEN_4412 : _GEN_4403; // @[NulCtrlMP.scala 789:23]
  wire  _GEN_4422 = cnt[20] ? _GEN_4413 : _GEN_4404; // @[NulCtrlMP.scala 789:23]
  wire  _GEN_4423 = cnt[20] ? _GEN_4414 : _GEN_4405; // @[NulCtrlMP.scala 789:23]
  wire [31:0] _GEN_4424 = cnt[20] ? _GEN_4415 : _GEN_4406; // @[NulCtrlMP.scala 789:23]
  wire [31:0] _GEN_4425 = cnt[20] ? _GEN_4416 : _GEN_4407; // @[NulCtrlMP.scala 789:23]
  wire [31:0] _GEN_4426 = cnt[20] ? _GEN_4417 : _GEN_4408; // @[NulCtrlMP.scala 789:23]
  wire [31:0] _GEN_4427 = cnt[20] ? _GEN_4418 : _GEN_4409; // @[NulCtrlMP.scala 789:23]
  wire [128:0] _GEN_4428 = cnt[20] ? _GEN_4419 : _GEN_4410; // @[NulCtrlMP.scala 789:23]
  wire  _GEN_4429 = _GEN_145 | _GEN_4420; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4430 = _GEN_146 | _GEN_4421; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4431 = _GEN_147 | _GEN_4422; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4432 = _GEN_148 | _GEN_4423; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4433 = 2'h0 == opidx ? 32'h773423 : _GEN_4424; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4434 = 2'h1 == opidx ? 32'h773423 : _GEN_4425; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4435 = 2'h2 == opidx ? 32'h773423 : _GEN_4426; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4436 = 2'h3 == opidx ? 32'h773423 : _GEN_4427; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4437 = _GEN_1180 ? _cnt_T : _GEN_4428; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4438 = cnt[21] ? _GEN_4429 : _GEN_4420; // @[NulCtrlMP.scala 790:23]
  wire  _GEN_4439 = cnt[21] ? _GEN_4430 : _GEN_4421; // @[NulCtrlMP.scala 790:23]
  wire  _GEN_4440 = cnt[21] ? _GEN_4431 : _GEN_4422; // @[NulCtrlMP.scala 790:23]
  wire  _GEN_4441 = cnt[21] ? _GEN_4432 : _GEN_4423; // @[NulCtrlMP.scala 790:23]
  wire [31:0] _GEN_4442 = cnt[21] ? _GEN_4433 : _GEN_4424; // @[NulCtrlMP.scala 790:23]
  wire [31:0] _GEN_4443 = cnt[21] ? _GEN_4434 : _GEN_4425; // @[NulCtrlMP.scala 790:23]
  wire [31:0] _GEN_4444 = cnt[21] ? _GEN_4435 : _GEN_4426; // @[NulCtrlMP.scala 790:23]
  wire [31:0] _GEN_4445 = cnt[21] ? _GEN_4436 : _GEN_4427; // @[NulCtrlMP.scala 790:23]
  wire [128:0] _GEN_4446 = cnt[21] ? _GEN_4437 : _GEN_4428; // @[NulCtrlMP.scala 790:23]
  wire  _GEN_4447 = _GEN_145 | _GEN_4438; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4448 = _GEN_146 | _GEN_4439; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4449 = _GEN_147 | _GEN_4440; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4450 = _GEN_148 | _GEN_4441; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4451 = 2'h0 == opidx ? 32'h873823 : _GEN_4442; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4452 = 2'h1 == opidx ? 32'h873823 : _GEN_4443; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4453 = 2'h2 == opidx ? 32'h873823 : _GEN_4444; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4454 = 2'h3 == opidx ? 32'h873823 : _GEN_4445; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4455 = _GEN_1180 ? _cnt_T : _GEN_4446; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4456 = cnt[22] ? _GEN_4447 : _GEN_4438; // @[NulCtrlMP.scala 791:23]
  wire  _GEN_4457 = cnt[22] ? _GEN_4448 : _GEN_4439; // @[NulCtrlMP.scala 791:23]
  wire  _GEN_4458 = cnt[22] ? _GEN_4449 : _GEN_4440; // @[NulCtrlMP.scala 791:23]
  wire  _GEN_4459 = cnt[22] ? _GEN_4450 : _GEN_4441; // @[NulCtrlMP.scala 791:23]
  wire [31:0] _GEN_4460 = cnt[22] ? _GEN_4451 : _GEN_4442; // @[NulCtrlMP.scala 791:23]
  wire [31:0] _GEN_4461 = cnt[22] ? _GEN_4452 : _GEN_4443; // @[NulCtrlMP.scala 791:23]
  wire [31:0] _GEN_4462 = cnt[22] ? _GEN_4453 : _GEN_4444; // @[NulCtrlMP.scala 791:23]
  wire [31:0] _GEN_4463 = cnt[22] ? _GEN_4454 : _GEN_4445; // @[NulCtrlMP.scala 791:23]
  wire [128:0] _GEN_4464 = cnt[22] ? _GEN_4455 : _GEN_4446; // @[NulCtrlMP.scala 791:23]
  wire  _GEN_4465 = _GEN_145 | _GEN_4456; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4466 = _GEN_146 | _GEN_4457; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4467 = _GEN_147 | _GEN_4458; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4468 = _GEN_148 | _GEN_4459; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4469 = 2'h0 == opidx ? 32'h973c23 : _GEN_4460; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4470 = 2'h1 == opidx ? 32'h973c23 : _GEN_4461; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4471 = 2'h2 == opidx ? 32'h973c23 : _GEN_4462; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4472 = 2'h3 == opidx ? 32'h973c23 : _GEN_4463; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4473 = _GEN_1180 ? _cnt_T : _GEN_4464; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4474 = cnt[23] ? _GEN_4465 : _GEN_4456; // @[NulCtrlMP.scala 792:23]
  wire  _GEN_4475 = cnt[23] ? _GEN_4466 : _GEN_4457; // @[NulCtrlMP.scala 792:23]
  wire  _GEN_4476 = cnt[23] ? _GEN_4467 : _GEN_4458; // @[NulCtrlMP.scala 792:23]
  wire  _GEN_4477 = cnt[23] ? _GEN_4468 : _GEN_4459; // @[NulCtrlMP.scala 792:23]
  wire [31:0] _GEN_4478 = cnt[23] ? _GEN_4469 : _GEN_4460; // @[NulCtrlMP.scala 792:23]
  wire [31:0] _GEN_4479 = cnt[23] ? _GEN_4470 : _GEN_4461; // @[NulCtrlMP.scala 792:23]
  wire [31:0] _GEN_4480 = cnt[23] ? _GEN_4471 : _GEN_4462; // @[NulCtrlMP.scala 792:23]
  wire [31:0] _GEN_4481 = cnt[23] ? _GEN_4472 : _GEN_4463; // @[NulCtrlMP.scala 792:23]
  wire [128:0] _GEN_4482 = cnt[23] ? _GEN_4473 : _GEN_4464; // @[NulCtrlMP.scala 792:23]
  wire  _GEN_4483 = _GEN_145 | _GEN_4474; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4484 = _GEN_146 | _GEN_4475; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4485 = _GEN_147 | _GEN_4476; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4486 = _GEN_148 | _GEN_4477; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4487 = 2'h0 == opidx ? 32'h2a73023 : _GEN_4478; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4488 = 2'h1 == opidx ? 32'h2a73023 : _GEN_4479; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4489 = 2'h2 == opidx ? 32'h2a73023 : _GEN_4480; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4490 = 2'h3 == opidx ? 32'h2a73023 : _GEN_4481; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4491 = _GEN_1180 ? _cnt_T : _GEN_4482; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4492 = cnt[24] ? _GEN_4483 : _GEN_4474; // @[NulCtrlMP.scala 793:23]
  wire  _GEN_4493 = cnt[24] ? _GEN_4484 : _GEN_4475; // @[NulCtrlMP.scala 793:23]
  wire  _GEN_4494 = cnt[24] ? _GEN_4485 : _GEN_4476; // @[NulCtrlMP.scala 793:23]
  wire  _GEN_4495 = cnt[24] ? _GEN_4486 : _GEN_4477; // @[NulCtrlMP.scala 793:23]
  wire [31:0] _GEN_4496 = cnt[24] ? _GEN_4487 : _GEN_4478; // @[NulCtrlMP.scala 793:23]
  wire [31:0] _GEN_4497 = cnt[24] ? _GEN_4488 : _GEN_4479; // @[NulCtrlMP.scala 793:23]
  wire [31:0] _GEN_4498 = cnt[24] ? _GEN_4489 : _GEN_4480; // @[NulCtrlMP.scala 793:23]
  wire [31:0] _GEN_4499 = cnt[24] ? _GEN_4490 : _GEN_4481; // @[NulCtrlMP.scala 793:23]
  wire [128:0] _GEN_4500 = cnt[24] ? _GEN_4491 : _GEN_4482; // @[NulCtrlMP.scala 793:23]
  wire  _GEN_4501 = _GEN_145 | _GEN_4492; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4502 = _GEN_146 | _GEN_4493; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4503 = _GEN_147 | _GEN_4494; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4504 = _GEN_148 | _GEN_4495; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4505 = 2'h0 == opidx ? 32'h2b73423 : _GEN_4496; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4506 = 2'h1 == opidx ? 32'h2b73423 : _GEN_4497; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4507 = 2'h2 == opidx ? 32'h2b73423 : _GEN_4498; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4508 = 2'h3 == opidx ? 32'h2b73423 : _GEN_4499; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4509 = _GEN_1180 ? _cnt_T : _GEN_4500; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4510 = cnt[25] ? _GEN_4501 : _GEN_4492; // @[NulCtrlMP.scala 794:23]
  wire  _GEN_4511 = cnt[25] ? _GEN_4502 : _GEN_4493; // @[NulCtrlMP.scala 794:23]
  wire  _GEN_4512 = cnt[25] ? _GEN_4503 : _GEN_4494; // @[NulCtrlMP.scala 794:23]
  wire  _GEN_4513 = cnt[25] ? _GEN_4504 : _GEN_4495; // @[NulCtrlMP.scala 794:23]
  wire [31:0] _GEN_4514 = cnt[25] ? _GEN_4505 : _GEN_4496; // @[NulCtrlMP.scala 794:23]
  wire [31:0] _GEN_4515 = cnt[25] ? _GEN_4506 : _GEN_4497; // @[NulCtrlMP.scala 794:23]
  wire [31:0] _GEN_4516 = cnt[25] ? _GEN_4507 : _GEN_4498; // @[NulCtrlMP.scala 794:23]
  wire [31:0] _GEN_4517 = cnt[25] ? _GEN_4508 : _GEN_4499; // @[NulCtrlMP.scala 794:23]
  wire [128:0] _GEN_4518 = cnt[25] ? _GEN_4509 : _GEN_4500; // @[NulCtrlMP.scala 794:23]
  wire  _GEN_4519 = _GEN_145 | _GEN_4510; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4520 = _GEN_146 | _GEN_4511; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4521 = _GEN_147 | _GEN_4512; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4522 = _GEN_148 | _GEN_4513; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4523 = 2'h0 == opidx ? 32'h2c73823 : _GEN_4514; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4524 = 2'h1 == opidx ? 32'h2c73823 : _GEN_4515; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4525 = 2'h2 == opidx ? 32'h2c73823 : _GEN_4516; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4526 = 2'h3 == opidx ? 32'h2c73823 : _GEN_4517; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4527 = _GEN_1180 ? _cnt_T : _GEN_4518; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4528 = cnt[26] ? _GEN_4519 : _GEN_4510; // @[NulCtrlMP.scala 795:23]
  wire  _GEN_4529 = cnt[26] ? _GEN_4520 : _GEN_4511; // @[NulCtrlMP.scala 795:23]
  wire  _GEN_4530 = cnt[26] ? _GEN_4521 : _GEN_4512; // @[NulCtrlMP.scala 795:23]
  wire  _GEN_4531 = cnt[26] ? _GEN_4522 : _GEN_4513; // @[NulCtrlMP.scala 795:23]
  wire [31:0] _GEN_4532 = cnt[26] ? _GEN_4523 : _GEN_4514; // @[NulCtrlMP.scala 795:23]
  wire [31:0] _GEN_4533 = cnt[26] ? _GEN_4524 : _GEN_4515; // @[NulCtrlMP.scala 795:23]
  wire [31:0] _GEN_4534 = cnt[26] ? _GEN_4525 : _GEN_4516; // @[NulCtrlMP.scala 795:23]
  wire [31:0] _GEN_4535 = cnt[26] ? _GEN_4526 : _GEN_4517; // @[NulCtrlMP.scala 795:23]
  wire [128:0] _GEN_4536 = cnt[26] ? _GEN_4527 : _GEN_4518; // @[NulCtrlMP.scala 795:23]
  wire  _GEN_4537 = _GEN_145 | _GEN_4528; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4538 = _GEN_146 | _GEN_4529; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4539 = _GEN_147 | _GEN_4530; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4540 = _GEN_148 | _GEN_4531; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4541 = 2'h0 == opidx ? 32'h2d73c23 : _GEN_4532; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4542 = 2'h1 == opidx ? 32'h2d73c23 : _GEN_4533; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4543 = 2'h2 == opidx ? 32'h2d73c23 : _GEN_4534; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4544 = 2'h3 == opidx ? 32'h2d73c23 : _GEN_4535; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4545 = _GEN_1180 ? _cnt_T : _GEN_4536; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4546 = cnt[27] ? _GEN_4537 : _GEN_4528; // @[NulCtrlMP.scala 796:23]
  wire  _GEN_4547 = cnt[27] ? _GEN_4538 : _GEN_4529; // @[NulCtrlMP.scala 796:23]
  wire  _GEN_4548 = cnt[27] ? _GEN_4539 : _GEN_4530; // @[NulCtrlMP.scala 796:23]
  wire  _GEN_4549 = cnt[27] ? _GEN_4540 : _GEN_4531; // @[NulCtrlMP.scala 796:23]
  wire [31:0] _GEN_4550 = cnt[27] ? _GEN_4541 : _GEN_4532; // @[NulCtrlMP.scala 796:23]
  wire [31:0] _GEN_4551 = cnt[27] ? _GEN_4542 : _GEN_4533; // @[NulCtrlMP.scala 796:23]
  wire [31:0] _GEN_4552 = cnt[27] ? _GEN_4543 : _GEN_4534; // @[NulCtrlMP.scala 796:23]
  wire [31:0] _GEN_4553 = cnt[27] ? _GEN_4544 : _GEN_4535; // @[NulCtrlMP.scala 796:23]
  wire [128:0] _GEN_4554 = cnt[27] ? _GEN_4545 : _GEN_4536; // @[NulCtrlMP.scala 796:23]
  wire  _GEN_4555 = _GEN_145 | _GEN_4546; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4556 = _GEN_146 | _GEN_4547; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4557 = _GEN_147 | _GEN_4548; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4558 = _GEN_148 | _GEN_4549; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4559 = 2'h0 == opidx ? 32'h4028293 : _GEN_4550; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4560 = 2'h1 == opidx ? 32'h4028293 : _GEN_4551; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4561 = 2'h2 == opidx ? 32'h4028293 : _GEN_4552; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4562 = 2'h3 == opidx ? 32'h4028293 : _GEN_4553; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4563 = _GEN_1180 ? _cnt_T : _GEN_4554; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4564 = cnt[28] ? _GEN_4555 : _GEN_4546; // @[NulCtrlMP.scala 797:23]
  wire  _GEN_4565 = cnt[28] ? _GEN_4556 : _GEN_4547; // @[NulCtrlMP.scala 797:23]
  wire  _GEN_4566 = cnt[28] ? _GEN_4557 : _GEN_4548; // @[NulCtrlMP.scala 797:23]
  wire  _GEN_4567 = cnt[28] ? _GEN_4558 : _GEN_4549; // @[NulCtrlMP.scala 797:23]
  wire [31:0] _GEN_4568 = cnt[28] ? _GEN_4559 : _GEN_4550; // @[NulCtrlMP.scala 797:23]
  wire [31:0] _GEN_4569 = cnt[28] ? _GEN_4560 : _GEN_4551; // @[NulCtrlMP.scala 797:23]
  wire [31:0] _GEN_4570 = cnt[28] ? _GEN_4561 : _GEN_4552; // @[NulCtrlMP.scala 797:23]
  wire [31:0] _GEN_4571 = cnt[28] ? _GEN_4562 : _GEN_4553; // @[NulCtrlMP.scala 797:23]
  wire [128:0] _GEN_4572 = cnt[28] ? _GEN_4563 : _GEN_4554; // @[NulCtrlMP.scala 797:23]
  wire  _GEN_4573 = _GEN_145 | _GEN_4564; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4574 = _GEN_146 | _GEN_4565; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4575 = _GEN_147 | _GEN_4566; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4576 = _GEN_148 | _GEN_4567; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4577 = 2'h0 == opidx ? 32'h4070713 : _GEN_4568; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4578 = 2'h1 == opidx ? 32'h4070713 : _GEN_4569; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4579 = 2'h2 == opidx ? 32'h4070713 : _GEN_4570; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4580 = 2'h3 == opidx ? 32'h4070713 : _GEN_4571; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4581 = _GEN_1180 ? _cnt_T : _GEN_4572; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4582 = cnt[29] ? _GEN_4573 : _GEN_4564; // @[NulCtrlMP.scala 798:23]
  wire  _GEN_4583 = cnt[29] ? _GEN_4574 : _GEN_4565; // @[NulCtrlMP.scala 798:23]
  wire  _GEN_4584 = cnt[29] ? _GEN_4575 : _GEN_4566; // @[NulCtrlMP.scala 798:23]
  wire  _GEN_4585 = cnt[29] ? _GEN_4576 : _GEN_4567; // @[NulCtrlMP.scala 798:23]
  wire [31:0] _GEN_4586 = cnt[29] ? _GEN_4577 : _GEN_4568; // @[NulCtrlMP.scala 798:23]
  wire [31:0] _GEN_4587 = cnt[29] ? _GEN_4578 : _GEN_4569; // @[NulCtrlMP.scala 798:23]
  wire [31:0] _GEN_4588 = cnt[29] ? _GEN_4579 : _GEN_4570; // @[NulCtrlMP.scala 798:23]
  wire [31:0] _GEN_4589 = cnt[29] ? _GEN_4580 : _GEN_4571; // @[NulCtrlMP.scala 798:23]
  wire [128:0] _GEN_4590 = cnt[29] ? _GEN_4581 : _GEN_4572; // @[NulCtrlMP.scala 798:23]
  wire  _GEN_4591 = _GEN_145 | _GEN_4009; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_4592 = _GEN_146 | _GEN_4010; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_4593 = _GEN_147 | _GEN_4011; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_4594 = _GEN_148 | _GEN_4012; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_4595 = ~_GEN_1252 ? _cnt_T : _GEN_4590; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_4596 = cnt[30] ? _GEN_4591 : _GEN_4009; // @[NulCtrlMP.scala 799:23]
  wire  _GEN_4597 = cnt[30] ? _GEN_4592 : _GEN_4010; // @[NulCtrlMP.scala 799:23]
  wire  _GEN_4598 = cnt[30] ? _GEN_4593 : _GEN_4011; // @[NulCtrlMP.scala 799:23]
  wire  _GEN_4599 = cnt[30] ? _GEN_4594 : _GEN_4012; // @[NulCtrlMP.scala 799:23]
  wire [128:0] _GEN_4600 = cnt[30] ? _GEN_4595 : _GEN_4590; // @[NulCtrlMP.scala 799:23]
  wire [128:0] _GEN_4601 = pg_loop_cnt < 8'h3f ? 129'h1000 : _cnt_T; // @[NulCtrlMP.scala 801:38 802:21 805:21]
  wire [128:0] _GEN_4603 = cnt[31] ? _GEN_4601 : _GEN_4600; // @[NulCtrlMP.scala 800:23]
  wire  _GEN_4605 = _GEN_145 | _GEN_4582; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4606 = _GEN_146 | _GEN_4583; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4607 = _GEN_147 | _GEN_4584; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_4608 = _GEN_148 | _GEN_4585; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_4609 = 2'h0 == opidx ? 32'h330000f : _GEN_4586; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4610 = 2'h1 == opidx ? 32'h330000f : _GEN_4587; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4611 = 2'h2 == opidx ? 32'h330000f : _GEN_4588; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_4612 = 2'h3 == opidx ? 32'h330000f : _GEN_4589; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_4613 = _GEN_1180 ? _cnt_T : _GEN_4603; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_4614 = cnt[32] ? _GEN_4605 : _GEN_4582; // @[NulCtrlMP.scala 809:23]
  wire  _GEN_4615 = cnt[32] ? _GEN_4606 : _GEN_4583; // @[NulCtrlMP.scala 809:23]
  wire  _GEN_4616 = cnt[32] ? _GEN_4607 : _GEN_4584; // @[NulCtrlMP.scala 809:23]
  wire  _GEN_4617 = cnt[32] ? _GEN_4608 : _GEN_4585; // @[NulCtrlMP.scala 809:23]
  wire [31:0] _GEN_4618 = cnt[32] ? _GEN_4609 : _GEN_4586; // @[NulCtrlMP.scala 809:23]
  wire [31:0] _GEN_4619 = cnt[32] ? _GEN_4610 : _GEN_4587; // @[NulCtrlMP.scala 809:23]
  wire [31:0] _GEN_4620 = cnt[32] ? _GEN_4611 : _GEN_4588; // @[NulCtrlMP.scala 809:23]
  wire [31:0] _GEN_4621 = cnt[32] ? _GEN_4612 : _GEN_4589; // @[NulCtrlMP.scala 809:23]
  wire [128:0] _GEN_4622 = cnt[32] ? _GEN_4613 : _GEN_4603; // @[NulCtrlMP.scala 809:23]
  wire  _GEN_4623 = _GEN_145 | _GEN_4596; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_4624 = _GEN_146 | _GEN_4597; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_4625 = _GEN_147 | _GEN_4598; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_4626 = _GEN_148 | _GEN_4599; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_4627 = ~_GEN_1252 ? _cnt_T : _GEN_4622; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_4628 = cnt[33] ? _GEN_4623 : _GEN_4596; // @[NulCtrlMP.scala 810:23]
  wire  _GEN_4629 = cnt[33] ? _GEN_4624 : _GEN_4597; // @[NulCtrlMP.scala 810:23]
  wire  _GEN_4630 = cnt[33] ? _GEN_4625 : _GEN_4598; // @[NulCtrlMP.scala 810:23]
  wire  _GEN_4631 = cnt[33] ? _GEN_4626 : _GEN_4599; // @[NulCtrlMP.scala 810:23]
  wire [128:0] _GEN_4632 = cnt[33] ? _GEN_4627 : _GEN_4622; // @[NulCtrlMP.scala 810:23]
  wire  _GEN_4633 = _GEN_145 | _GEN_4254; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4634 = _GEN_146 | _GEN_4255; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4635 = _GEN_147 | _GEN_4256; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4636 = _GEN_148 | _GEN_4257; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4637 = 2'h0 == opidx ? 5'h5 : _GEN_4258; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4638 = 2'h1 == opidx ? 5'h5 : _GEN_4259; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4639 = 2'h2 == opidx ? 5'h5 : _GEN_4260; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4640 = 2'h3 == opidx ? 5'h5 : _GEN_4261; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4641 = 2'h0 == opidx ? regback_0 : _GEN_4262; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4642 = 2'h1 == opidx ? regback_0 : _GEN_4263; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4643 = 2'h2 == opidx ? regback_0 : _GEN_4264; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4644 = 2'h3 == opidx ? regback_0 : _GEN_4265; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4645 = ~_GEN_1128 ? _cnt_T : _GEN_4632; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4646 = cnt[34] ? _GEN_4633 : _GEN_4254; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4647 = cnt[34] ? _GEN_4634 : _GEN_4255; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4648 = cnt[34] ? _GEN_4635 : _GEN_4256; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4649 = cnt[34] ? _GEN_4636 : _GEN_4257; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4650 = cnt[34] ? _GEN_4637 : _GEN_4258; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4651 = cnt[34] ? _GEN_4638 : _GEN_4259; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4652 = cnt[34] ? _GEN_4639 : _GEN_4260; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4653 = cnt[34] ? _GEN_4640 : _GEN_4261; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4654 = cnt[34] ? _GEN_4641 : _GEN_4262; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4655 = cnt[34] ? _GEN_4642 : _GEN_4263; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4656 = cnt[34] ? _GEN_4643 : _GEN_4264; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4657 = cnt[34] ? _GEN_4644 : _GEN_4265; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4658 = cnt[34] ? _GEN_4645 : _GEN_4632; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4659 = _GEN_145 | _GEN_4646; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4660 = _GEN_146 | _GEN_4647; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4661 = _GEN_147 | _GEN_4648; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4662 = _GEN_148 | _GEN_4649; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4663 = 2'h0 == opidx ? 5'h6 : _GEN_4650; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4664 = 2'h1 == opidx ? 5'h6 : _GEN_4651; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4665 = 2'h2 == opidx ? 5'h6 : _GEN_4652; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4666 = 2'h3 == opidx ? 5'h6 : _GEN_4653; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4667 = 2'h0 == opidx ? regback_1 : _GEN_4654; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4668 = 2'h1 == opidx ? regback_1 : _GEN_4655; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4669 = 2'h2 == opidx ? regback_1 : _GEN_4656; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4670 = 2'h3 == opidx ? regback_1 : _GEN_4657; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4671 = ~_GEN_1128 ? _cnt_T : _GEN_4658; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4672 = cnt[35] ? _GEN_4659 : _GEN_4646; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4673 = cnt[35] ? _GEN_4660 : _GEN_4647; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4674 = cnt[35] ? _GEN_4661 : _GEN_4648; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4675 = cnt[35] ? _GEN_4662 : _GEN_4649; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4676 = cnt[35] ? _GEN_4663 : _GEN_4650; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4677 = cnt[35] ? _GEN_4664 : _GEN_4651; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4678 = cnt[35] ? _GEN_4665 : _GEN_4652; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4679 = cnt[35] ? _GEN_4666 : _GEN_4653; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4680 = cnt[35] ? _GEN_4667 : _GEN_4654; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4681 = cnt[35] ? _GEN_4668 : _GEN_4655; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4682 = cnt[35] ? _GEN_4669 : _GEN_4656; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4683 = cnt[35] ? _GEN_4670 : _GEN_4657; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4684 = cnt[35] ? _GEN_4671 : _GEN_4658; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4685 = _GEN_145 | _GEN_4672; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4686 = _GEN_146 | _GEN_4673; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4687 = _GEN_147 | _GEN_4674; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4688 = _GEN_148 | _GEN_4675; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4689 = 2'h0 == opidx ? 5'h7 : _GEN_4676; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4690 = 2'h1 == opidx ? 5'h7 : _GEN_4677; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4691 = 2'h2 == opidx ? 5'h7 : _GEN_4678; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4692 = 2'h3 == opidx ? 5'h7 : _GEN_4679; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4693 = 2'h0 == opidx ? regback_2 : _GEN_4680; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4694 = 2'h1 == opidx ? regback_2 : _GEN_4681; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4695 = 2'h2 == opidx ? regback_2 : _GEN_4682; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4696 = 2'h3 == opidx ? regback_2 : _GEN_4683; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4697 = ~_GEN_1128 ? _cnt_T : _GEN_4684; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4698 = cnt[36] ? _GEN_4685 : _GEN_4672; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4699 = cnt[36] ? _GEN_4686 : _GEN_4673; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4700 = cnt[36] ? _GEN_4687 : _GEN_4674; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4701 = cnt[36] ? _GEN_4688 : _GEN_4675; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4702 = cnt[36] ? _GEN_4689 : _GEN_4676; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4703 = cnt[36] ? _GEN_4690 : _GEN_4677; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4704 = cnt[36] ? _GEN_4691 : _GEN_4678; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4705 = cnt[36] ? _GEN_4692 : _GEN_4679; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4706 = cnt[36] ? _GEN_4693 : _GEN_4680; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4707 = cnt[36] ? _GEN_4694 : _GEN_4681; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4708 = cnt[36] ? _GEN_4695 : _GEN_4682; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4709 = cnt[36] ? _GEN_4696 : _GEN_4683; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4710 = cnt[36] ? _GEN_4697 : _GEN_4684; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4711 = _GEN_145 | _GEN_4698; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4712 = _GEN_146 | _GEN_4699; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4713 = _GEN_147 | _GEN_4700; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4714 = _GEN_148 | _GEN_4701; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4715 = 2'h0 == opidx ? 5'h8 : _GEN_4702; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4716 = 2'h1 == opidx ? 5'h8 : _GEN_4703; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4717 = 2'h2 == opidx ? 5'h8 : _GEN_4704; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4718 = 2'h3 == opidx ? 5'h8 : _GEN_4705; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4719 = 2'h0 == opidx ? regback_3 : _GEN_4706; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4720 = 2'h1 == opidx ? regback_3 : _GEN_4707; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4721 = 2'h2 == opidx ? regback_3 : _GEN_4708; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4722 = 2'h3 == opidx ? regback_3 : _GEN_4709; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4723 = ~_GEN_1128 ? _cnt_T : _GEN_4710; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4724 = cnt[37] ? _GEN_4711 : _GEN_4698; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4725 = cnt[37] ? _GEN_4712 : _GEN_4699; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4726 = cnt[37] ? _GEN_4713 : _GEN_4700; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4727 = cnt[37] ? _GEN_4714 : _GEN_4701; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4728 = cnt[37] ? _GEN_4715 : _GEN_4702; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4729 = cnt[37] ? _GEN_4716 : _GEN_4703; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4730 = cnt[37] ? _GEN_4717 : _GEN_4704; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4731 = cnt[37] ? _GEN_4718 : _GEN_4705; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4732 = cnt[37] ? _GEN_4719 : _GEN_4706; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4733 = cnt[37] ? _GEN_4720 : _GEN_4707; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4734 = cnt[37] ? _GEN_4721 : _GEN_4708; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4735 = cnt[37] ? _GEN_4722 : _GEN_4709; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4736 = cnt[37] ? _GEN_4723 : _GEN_4710; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4737 = _GEN_145 | _GEN_4724; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4738 = _GEN_146 | _GEN_4725; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4739 = _GEN_147 | _GEN_4726; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4740 = _GEN_148 | _GEN_4727; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4741 = 2'h0 == opidx ? 5'h9 : _GEN_4728; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4742 = 2'h1 == opidx ? 5'h9 : _GEN_4729; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4743 = 2'h2 == opidx ? 5'h9 : _GEN_4730; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4744 = 2'h3 == opidx ? 5'h9 : _GEN_4731; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4745 = 2'h0 == opidx ? regback_4 : _GEN_4732; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4746 = 2'h1 == opidx ? regback_4 : _GEN_4733; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4747 = 2'h2 == opidx ? regback_4 : _GEN_4734; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4748 = 2'h3 == opidx ? regback_4 : _GEN_4735; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4749 = ~_GEN_1128 ? _cnt_T : _GEN_4736; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4750 = cnt[38] ? _GEN_4737 : _GEN_4724; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4751 = cnt[38] ? _GEN_4738 : _GEN_4725; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4752 = cnt[38] ? _GEN_4739 : _GEN_4726; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4753 = cnt[38] ? _GEN_4740 : _GEN_4727; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4754 = cnt[38] ? _GEN_4741 : _GEN_4728; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4755 = cnt[38] ? _GEN_4742 : _GEN_4729; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4756 = cnt[38] ? _GEN_4743 : _GEN_4730; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4757 = cnt[38] ? _GEN_4744 : _GEN_4731; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4758 = cnt[38] ? _GEN_4745 : _GEN_4732; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4759 = cnt[38] ? _GEN_4746 : _GEN_4733; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4760 = cnt[38] ? _GEN_4747 : _GEN_4734; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4761 = cnt[38] ? _GEN_4748 : _GEN_4735; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4762 = cnt[38] ? _GEN_4749 : _GEN_4736; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4763 = _GEN_145 | _GEN_4750; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4764 = _GEN_146 | _GEN_4751; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4765 = _GEN_147 | _GEN_4752; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4766 = _GEN_148 | _GEN_4753; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4767 = 2'h0 == opidx ? 5'ha : _GEN_4754; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4768 = 2'h1 == opidx ? 5'ha : _GEN_4755; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4769 = 2'h2 == opidx ? 5'ha : _GEN_4756; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4770 = 2'h3 == opidx ? 5'ha : _GEN_4757; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4771 = 2'h0 == opidx ? regback_5 : _GEN_4758; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4772 = 2'h1 == opidx ? regback_5 : _GEN_4759; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4773 = 2'h2 == opidx ? regback_5 : _GEN_4760; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4774 = 2'h3 == opidx ? regback_5 : _GEN_4761; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4775 = ~_GEN_1128 ? _cnt_T : _GEN_4762; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4776 = cnt[39] ? _GEN_4763 : _GEN_4750; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4777 = cnt[39] ? _GEN_4764 : _GEN_4751; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4778 = cnt[39] ? _GEN_4765 : _GEN_4752; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4779 = cnt[39] ? _GEN_4766 : _GEN_4753; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4780 = cnt[39] ? _GEN_4767 : _GEN_4754; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4781 = cnt[39] ? _GEN_4768 : _GEN_4755; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4782 = cnt[39] ? _GEN_4769 : _GEN_4756; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4783 = cnt[39] ? _GEN_4770 : _GEN_4757; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4784 = cnt[39] ? _GEN_4771 : _GEN_4758; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4785 = cnt[39] ? _GEN_4772 : _GEN_4759; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4786 = cnt[39] ? _GEN_4773 : _GEN_4760; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4787 = cnt[39] ? _GEN_4774 : _GEN_4761; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4788 = cnt[39] ? _GEN_4775 : _GEN_4762; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4789 = _GEN_145 | _GEN_4776; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4790 = _GEN_146 | _GEN_4777; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4791 = _GEN_147 | _GEN_4778; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4792 = _GEN_148 | _GEN_4779; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4793 = 2'h0 == opidx ? 5'hb : _GEN_4780; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4794 = 2'h1 == opidx ? 5'hb : _GEN_4781; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4795 = 2'h2 == opidx ? 5'hb : _GEN_4782; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4796 = 2'h3 == opidx ? 5'hb : _GEN_4783; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4797 = 2'h0 == opidx ? regback_6 : _GEN_4784; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4798 = 2'h1 == opidx ? regback_6 : _GEN_4785; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4799 = 2'h2 == opidx ? regback_6 : _GEN_4786; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4800 = 2'h3 == opidx ? regback_6 : _GEN_4787; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4801 = ~_GEN_1128 ? _cnt_T : _GEN_4788; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4802 = cnt[40] ? _GEN_4789 : _GEN_4776; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4803 = cnt[40] ? _GEN_4790 : _GEN_4777; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4804 = cnt[40] ? _GEN_4791 : _GEN_4778; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4805 = cnt[40] ? _GEN_4792 : _GEN_4779; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4806 = cnt[40] ? _GEN_4793 : _GEN_4780; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4807 = cnt[40] ? _GEN_4794 : _GEN_4781; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4808 = cnt[40] ? _GEN_4795 : _GEN_4782; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4809 = cnt[40] ? _GEN_4796 : _GEN_4783; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4810 = cnt[40] ? _GEN_4797 : _GEN_4784; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4811 = cnt[40] ? _GEN_4798 : _GEN_4785; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4812 = cnt[40] ? _GEN_4799 : _GEN_4786; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4813 = cnt[40] ? _GEN_4800 : _GEN_4787; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4814 = cnt[40] ? _GEN_4801 : _GEN_4788; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4815 = _GEN_145 | _GEN_4802; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4816 = _GEN_146 | _GEN_4803; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4817 = _GEN_147 | _GEN_4804; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4818 = _GEN_148 | _GEN_4805; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4819 = 2'h0 == opidx ? 5'hc : _GEN_4806; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4820 = 2'h1 == opidx ? 5'hc : _GEN_4807; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4821 = 2'h2 == opidx ? 5'hc : _GEN_4808; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4822 = 2'h3 == opidx ? 5'hc : _GEN_4809; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4823 = 2'h0 == opidx ? regback_7 : _GEN_4810; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4824 = 2'h1 == opidx ? regback_7 : _GEN_4811; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4825 = 2'h2 == opidx ? regback_7 : _GEN_4812; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4826 = 2'h3 == opidx ? regback_7 : _GEN_4813; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4827 = ~_GEN_1128 ? _cnt_T : _GEN_4814; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4828 = cnt[41] ? _GEN_4815 : _GEN_4802; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4829 = cnt[41] ? _GEN_4816 : _GEN_4803; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4830 = cnt[41] ? _GEN_4817 : _GEN_4804; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4831 = cnt[41] ? _GEN_4818 : _GEN_4805; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4832 = cnt[41] ? _GEN_4819 : _GEN_4806; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4833 = cnt[41] ? _GEN_4820 : _GEN_4807; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4834 = cnt[41] ? _GEN_4821 : _GEN_4808; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4835 = cnt[41] ? _GEN_4822 : _GEN_4809; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4836 = cnt[41] ? _GEN_4823 : _GEN_4810; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4837 = cnt[41] ? _GEN_4824 : _GEN_4811; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4838 = cnt[41] ? _GEN_4825 : _GEN_4812; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4839 = cnt[41] ? _GEN_4826 : _GEN_4813; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4840 = cnt[41] ? _GEN_4827 : _GEN_4814; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4841 = _GEN_145 | _GEN_4828; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4842 = _GEN_146 | _GEN_4829; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4843 = _GEN_147 | _GEN_4830; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4844 = _GEN_148 | _GEN_4831; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4845 = 2'h0 == opidx ? 5'hd : _GEN_4832; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4846 = 2'h1 == opidx ? 5'hd : _GEN_4833; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4847 = 2'h2 == opidx ? 5'hd : _GEN_4834; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4848 = 2'h3 == opidx ? 5'hd : _GEN_4835; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4849 = 2'h0 == opidx ? regback_8 : _GEN_4836; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4850 = 2'h1 == opidx ? regback_8 : _GEN_4837; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4851 = 2'h2 == opidx ? regback_8 : _GEN_4838; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4852 = 2'h3 == opidx ? regback_8 : _GEN_4839; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4853 = ~_GEN_1128 ? _cnt_T : _GEN_4840; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4854 = cnt[42] ? _GEN_4841 : _GEN_4828; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4855 = cnt[42] ? _GEN_4842 : _GEN_4829; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4856 = cnt[42] ? _GEN_4843 : _GEN_4830; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4857 = cnt[42] ? _GEN_4844 : _GEN_4831; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4858 = cnt[42] ? _GEN_4845 : _GEN_4832; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4859 = cnt[42] ? _GEN_4846 : _GEN_4833; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4860 = cnt[42] ? _GEN_4847 : _GEN_4834; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4861 = cnt[42] ? _GEN_4848 : _GEN_4835; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4862 = cnt[42] ? _GEN_4849 : _GEN_4836; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4863 = cnt[42] ? _GEN_4850 : _GEN_4837; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4864 = cnt[42] ? _GEN_4851 : _GEN_4838; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4865 = cnt[42] ? _GEN_4852 : _GEN_4839; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4866 = cnt[42] ? _GEN_4853 : _GEN_4840; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4867 = _GEN_145 | _GEN_4854; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4868 = _GEN_146 | _GEN_4855; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4869 = _GEN_147 | _GEN_4856; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_4870 = _GEN_148 | _GEN_4857; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_4871 = 2'h0 == opidx ? 5'he : _GEN_4858; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4872 = 2'h1 == opidx ? 5'he : _GEN_4859; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4873 = 2'h2 == opidx ? 5'he : _GEN_4860; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_4874 = 2'h3 == opidx ? 5'he : _GEN_4861; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_4875 = 2'h0 == opidx ? regback_9 : _GEN_4862; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4876 = 2'h1 == opidx ? regback_9 : _GEN_4863; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4877 = 2'h2 == opidx ? regback_9 : _GEN_4864; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_4878 = 2'h3 == opidx ? regback_9 : _GEN_4865; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_4879 = ~_GEN_1128 ? _cnt_T : _GEN_4866; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_4880 = cnt[43] ? _GEN_4867 : _GEN_4854; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4881 = cnt[43] ? _GEN_4868 : _GEN_4855; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4882 = cnt[43] ? _GEN_4869 : _GEN_4856; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_4883 = cnt[43] ? _GEN_4870 : _GEN_4857; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4884 = cnt[43] ? _GEN_4871 : _GEN_4858; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4885 = cnt[43] ? _GEN_4872 : _GEN_4859; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4886 = cnt[43] ? _GEN_4873 : _GEN_4860; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_4887 = cnt[43] ? _GEN_4874 : _GEN_4861; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4888 = cnt[43] ? _GEN_4875 : _GEN_4862; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4889 = cnt[43] ? _GEN_4876 : _GEN_4863; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4890 = cnt[43] ? _GEN_4877 : _GEN_4864; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_4891 = cnt[43] ? _GEN_4878 : _GEN_4865; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4892 = cnt[43] ? _GEN_4879 : _GEN_4866; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_4893 = cnt[44] ? 129'h1 : _GEN_4892; // @[NulCtrlMP.scala 812:23 813:17]
  wire [4:0] _GEN_4894 = cnt[44] ? 5'h5 : _GEN_4014; // @[NulCtrlMP.scala 812:23 814:19]
  wire  _GEN_4895 = state == 5'h15 ? _GEN_4205 : _GEN_3982; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4896 = state == 5'h15 ? _GEN_4206 : _GEN_3983; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4897 = state == 5'h15 ? _GEN_4207 : _GEN_3984; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4898 = state == 5'h15 ? _GEN_4208 : _GEN_3985; // @[NulCtrlMP.scala 777:32]
  wire [4:0] _GEN_4899 = state == 5'h15 ? _GEN_4884 : _GEN_3986; // @[NulCtrlMP.scala 777:32]
  wire [4:0] _GEN_4900 = state == 5'h15 ? _GEN_4885 : _GEN_3987; // @[NulCtrlMP.scala 777:32]
  wire [4:0] _GEN_4901 = state == 5'h15 ? _GEN_4886 : _GEN_3988; // @[NulCtrlMP.scala 777:32]
  wire [4:0] _GEN_4902 = state == 5'h15 ? _GEN_4887 : _GEN_3989; // @[NulCtrlMP.scala 777:32]
  wire [128:0] _GEN_4903 = state == 5'h15 ? _GEN_4893 : _GEN_3990; // @[NulCtrlMP.scala 777:32]
  wire [63:0] _GEN_4904 = state == 5'h15 ? _GEN_4034 : _GEN_3991; // @[NulCtrlMP.scala 777:32]
  wire [63:0] _GEN_4905 = state == 5'h15 ? _GEN_4054 : _GEN_3992; // @[NulCtrlMP.scala 777:32]
  wire [63:0] _GEN_4906 = state == 5'h15 ? _GEN_4074 : _GEN_2439; // @[NulCtrlMP.scala 777:32]
  wire [63:0] _GEN_4907 = state == 5'h15 ? _GEN_4094 : regback_3; // @[NulCtrlMP.scala 346:26 777:32]
  wire [63:0] _GEN_4908 = state == 5'h15 ? _GEN_4114 : regback_4; // @[NulCtrlMP.scala 346:26 777:32]
  wire [63:0] _GEN_4909 = state == 5'h15 ? _GEN_4134 : regback_5; // @[NulCtrlMP.scala 346:26 777:32]
  wire [63:0] _GEN_4910 = state == 5'h15 ? _GEN_4154 : regback_6; // @[NulCtrlMP.scala 346:26 777:32]
  wire [63:0] _GEN_4911 = state == 5'h15 ? _GEN_4174 : regback_7; // @[NulCtrlMP.scala 346:26 777:32]
  wire [63:0] _GEN_4912 = state == 5'h15 ? _GEN_4194 : regback_8; // @[NulCtrlMP.scala 346:26 777:32]
  wire  _GEN_4914 = state == 5'h15 ? _GEN_4880 : _GEN_3993; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4915 = state == 5'h15 ? _GEN_4881 : _GEN_3994; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4916 = state == 5'h15 ? _GEN_4882 : _GEN_3995; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4917 = state == 5'h15 ? _GEN_4883 : _GEN_3996; // @[NulCtrlMP.scala 777:32]
  wire [63:0] _GEN_4918 = state == 5'h15 ? _GEN_4888 : _GEN_3997; // @[NulCtrlMP.scala 777:32]
  wire [63:0] _GEN_4919 = state == 5'h15 ? _GEN_4889 : _GEN_3998; // @[NulCtrlMP.scala 777:32]
  wire [63:0] _GEN_4920 = state == 5'h15 ? _GEN_4890 : _GEN_3999; // @[NulCtrlMP.scala 777:32]
  wire [63:0] _GEN_4921 = state == 5'h15 ? _GEN_4891 : _GEN_4000; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4922 = state == 5'h15 ? _GEN_4614 : _GEN_4001; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4923 = state == 5'h15 ? _GEN_4615 : _GEN_4002; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4924 = state == 5'h15 ? _GEN_4616 : _GEN_4003; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4925 = state == 5'h15 ? _GEN_4617 : _GEN_4004; // @[NulCtrlMP.scala 777:32]
  wire [31:0] _GEN_4926 = state == 5'h15 ? _GEN_4618 : _GEN_4005; // @[NulCtrlMP.scala 777:32]
  wire [31:0] _GEN_4927 = state == 5'h15 ? _GEN_4619 : _GEN_4006; // @[NulCtrlMP.scala 777:32]
  wire [31:0] _GEN_4928 = state == 5'h15 ? _GEN_4620 : _GEN_4007; // @[NulCtrlMP.scala 777:32]
  wire [31:0] _GEN_4929 = state == 5'h15 ? _GEN_4621 : _GEN_4008; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4930 = state == 5'h15 ? _GEN_4628 : _GEN_4009; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4931 = state == 5'h15 ? _GEN_4629 : _GEN_4010; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4932 = state == 5'h15 ? _GEN_4630 : _GEN_4011; // @[NulCtrlMP.scala 777:32]
  wire  _GEN_4933 = state == 5'h15 ? _GEN_4631 : _GEN_4012; // @[NulCtrlMP.scala 777:32]
  wire [4:0] _GEN_4935 = state == 5'h15 ? _GEN_4894 : _GEN_4014; // @[NulCtrlMP.scala 777:32]
  reg [63:0] pgbuf_div8_0; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_1; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_2; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_3; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_4; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_5; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_6; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_7; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_8; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_9; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_10; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_11; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_12; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_13; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_14; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_15; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_16; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_17; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_18; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_19; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_20; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_21; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_22; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_23; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_24; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_25; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_26; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_27; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_28; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_29; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_30; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_31; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_32; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_33; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_34; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_35; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_36; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_37; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_38; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_39; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_40; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_41; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_42; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_43; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_44; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_45; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_46; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_47; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_48; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_49; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_50; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_51; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_52; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_53; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_54; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_55; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_56; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_57; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_58; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_59; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_60; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_61; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_62; // @[NulCtrlMP.scala 818:29]
  reg [63:0] pgbuf_div8_63; // @[NulCtrlMP.scala 818:29]
  reg [11:0] pgbuf_uart_pos; // @[NulCtrlMP.scala 819:33]
  reg [11:0] pgbuf_cpu_pos; // @[NulCtrlMP.scala 820:32]
  wire  _GEN_4936 = _GEN_145 | _GEN_4895; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4937 = _GEN_146 | _GEN_4896; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4938 = _GEN_147 | _GEN_4897; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4939 = _GEN_148 | _GEN_4898; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4940 = 2'h0 == opidx ? 5'h5 : _GEN_4899; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4941 = 2'h1 == opidx ? 5'h5 : _GEN_4900; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4942 = 2'h2 == opidx ? 5'h5 : _GEN_4901; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4943 = 2'h3 == opidx ? 5'h5 : _GEN_4902; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4944 = _T_122 ? _cnt_T : _GEN_4903; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4945 = _T_122 ? _GEN_1349 : _GEN_4904; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_4946 = cnt[0] ? _GEN_4936 : _GEN_4895; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4947 = cnt[0] ? _GEN_4937 : _GEN_4896; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4948 = cnt[0] ? _GEN_4938 : _GEN_4897; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4949 = cnt[0] ? _GEN_4939 : _GEN_4898; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4950 = cnt[0] ? _GEN_4940 : _GEN_4899; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4951 = cnt[0] ? _GEN_4941 : _GEN_4900; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4952 = cnt[0] ? _GEN_4942 : _GEN_4901; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4953 = cnt[0] ? _GEN_4943 : _GEN_4902; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4954 = cnt[0] ? _GEN_4944 : _GEN_4903; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4955 = cnt[0] ? _GEN_4945 : _GEN_4904; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4956 = _GEN_145 | _GEN_4946; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4957 = _GEN_146 | _GEN_4947; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4958 = _GEN_147 | _GEN_4948; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4959 = _GEN_148 | _GEN_4949; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4960 = 2'h0 == opidx ? 5'h6 : _GEN_4950; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4961 = 2'h1 == opidx ? 5'h6 : _GEN_4951; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4962 = 2'h2 == opidx ? 5'h6 : _GEN_4952; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4963 = 2'h3 == opidx ? 5'h6 : _GEN_4953; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4964 = _T_122 ? _cnt_T : _GEN_4954; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4965 = _T_122 ? _GEN_1349 : _GEN_4905; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_4966 = cnt[1] ? _GEN_4956 : _GEN_4946; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4967 = cnt[1] ? _GEN_4957 : _GEN_4947; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4968 = cnt[1] ? _GEN_4958 : _GEN_4948; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4969 = cnt[1] ? _GEN_4959 : _GEN_4949; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4970 = cnt[1] ? _GEN_4960 : _GEN_4950; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4971 = cnt[1] ? _GEN_4961 : _GEN_4951; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4972 = cnt[1] ? _GEN_4962 : _GEN_4952; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4973 = cnt[1] ? _GEN_4963 : _GEN_4953; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4974 = cnt[1] ? _GEN_4964 : _GEN_4954; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4975 = cnt[1] ? _GEN_4965 : _GEN_4905; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4976 = _GEN_145 | _GEN_4966; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4977 = _GEN_146 | _GEN_4967; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4978 = _GEN_147 | _GEN_4968; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4979 = _GEN_148 | _GEN_4969; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_4980 = 2'h0 == opidx ? 5'h7 : _GEN_4970; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4981 = 2'h1 == opidx ? 5'h7 : _GEN_4971; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4982 = 2'h2 == opidx ? 5'h7 : _GEN_4972; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_4983 = 2'h3 == opidx ? 5'h7 : _GEN_4973; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_4984 = _T_122 ? _cnt_T : _GEN_4974; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_4985 = _T_122 ? _GEN_1349 : _GEN_4906; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_4986 = cnt[2] ? _GEN_4976 : _GEN_4966; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4987 = cnt[2] ? _GEN_4977 : _GEN_4967; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4988 = cnt[2] ? _GEN_4978 : _GEN_4968; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4989 = cnt[2] ? _GEN_4979 : _GEN_4969; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4990 = cnt[2] ? _GEN_4980 : _GEN_4970; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4991 = cnt[2] ? _GEN_4981 : _GEN_4971; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4992 = cnt[2] ? _GEN_4982 : _GEN_4972; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_4993 = cnt[2] ? _GEN_4983 : _GEN_4973; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_4994 = cnt[2] ? _GEN_4984 : _GEN_4974; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_4995 = cnt[2] ? _GEN_4985 : _GEN_4906; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_4996 = _GEN_145 | _GEN_4986; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4997 = _GEN_146 | _GEN_4987; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4998 = _GEN_147 | _GEN_4988; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_4999 = _GEN_148 | _GEN_4989; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5000 = 2'h0 == opidx ? 5'h8 : _GEN_4990; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5001 = 2'h1 == opidx ? 5'h8 : _GEN_4991; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5002 = 2'h2 == opidx ? 5'h8 : _GEN_4992; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5003 = 2'h3 == opidx ? 5'h8 : _GEN_4993; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_5004 = _T_122 ? _cnt_T : _GEN_4994; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_5005 = _T_122 ? _GEN_1349 : _GEN_4907; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_5006 = cnt[3] ? _GEN_4996 : _GEN_4986; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5007 = cnt[3] ? _GEN_4997 : _GEN_4987; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5008 = cnt[3] ? _GEN_4998 : _GEN_4988; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5009 = cnt[3] ? _GEN_4999 : _GEN_4989; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5010 = cnt[3] ? _GEN_5000 : _GEN_4990; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5011 = cnt[3] ? _GEN_5001 : _GEN_4991; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5012 = cnt[3] ? _GEN_5002 : _GEN_4992; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5013 = cnt[3] ? _GEN_5003 : _GEN_4993; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_5014 = cnt[3] ? _GEN_5004 : _GEN_4994; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_5015 = cnt[3] ? _GEN_5005 : _GEN_4907; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5016 = _GEN_145 | _GEN_5006; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5017 = _GEN_146 | _GEN_5007; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5018 = _GEN_147 | _GEN_5008; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5019 = _GEN_148 | _GEN_5009; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5020 = 2'h0 == opidx ? 5'h9 : _GEN_5010; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5021 = 2'h1 == opidx ? 5'h9 : _GEN_5011; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5022 = 2'h2 == opidx ? 5'h9 : _GEN_5012; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5023 = 2'h3 == opidx ? 5'h9 : _GEN_5013; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_5024 = _T_122 ? _cnt_T : _GEN_5014; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_5025 = _T_122 ? _GEN_1349 : _GEN_4908; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_5026 = cnt[4] ? _GEN_5016 : _GEN_5006; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5027 = cnt[4] ? _GEN_5017 : _GEN_5007; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5028 = cnt[4] ? _GEN_5018 : _GEN_5008; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5029 = cnt[4] ? _GEN_5019 : _GEN_5009; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5030 = cnt[4] ? _GEN_5020 : _GEN_5010; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5031 = cnt[4] ? _GEN_5021 : _GEN_5011; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5032 = cnt[4] ? _GEN_5022 : _GEN_5012; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5033 = cnt[4] ? _GEN_5023 : _GEN_5013; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_5034 = cnt[4] ? _GEN_5024 : _GEN_5014; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_5035 = cnt[4] ? _GEN_5025 : _GEN_4908; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5036 = _GEN_145 | _GEN_5026; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5037 = _GEN_146 | _GEN_5027; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5038 = _GEN_147 | _GEN_5028; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5039 = _GEN_148 | _GEN_5029; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5040 = 2'h0 == opidx ? 5'ha : _GEN_5030; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5041 = 2'h1 == opidx ? 5'ha : _GEN_5031; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5042 = 2'h2 == opidx ? 5'ha : _GEN_5032; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5043 = 2'h3 == opidx ? 5'ha : _GEN_5033; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_5044 = _T_122 ? _cnt_T : _GEN_5034; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_5045 = _T_122 ? _GEN_1349 : _GEN_4909; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_5046 = cnt[5] ? _GEN_5036 : _GEN_5026; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5047 = cnt[5] ? _GEN_5037 : _GEN_5027; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5048 = cnt[5] ? _GEN_5038 : _GEN_5028; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5049 = cnt[5] ? _GEN_5039 : _GEN_5029; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5050 = cnt[5] ? _GEN_5040 : _GEN_5030; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5051 = cnt[5] ? _GEN_5041 : _GEN_5031; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5052 = cnt[5] ? _GEN_5042 : _GEN_5032; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5053 = cnt[5] ? _GEN_5043 : _GEN_5033; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_5054 = cnt[5] ? _GEN_5044 : _GEN_5034; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_5055 = cnt[5] ? _GEN_5045 : _GEN_4909; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5056 = _GEN_145 | _GEN_5046; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5057 = _GEN_146 | _GEN_5047; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5058 = _GEN_147 | _GEN_5048; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5059 = _GEN_148 | _GEN_5049; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5060 = 2'h0 == opidx ? 5'hb : _GEN_5050; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5061 = 2'h1 == opidx ? 5'hb : _GEN_5051; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5062 = 2'h2 == opidx ? 5'hb : _GEN_5052; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5063 = 2'h3 == opidx ? 5'hb : _GEN_5053; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_5064 = _T_122 ? _cnt_T : _GEN_5054; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_5065 = _T_122 ? _GEN_1349 : _GEN_4910; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_5066 = cnt[6] ? _GEN_5056 : _GEN_5046; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5067 = cnt[6] ? _GEN_5057 : _GEN_5047; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5068 = cnt[6] ? _GEN_5058 : _GEN_5048; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5069 = cnt[6] ? _GEN_5059 : _GEN_5049; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5070 = cnt[6] ? _GEN_5060 : _GEN_5050; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5071 = cnt[6] ? _GEN_5061 : _GEN_5051; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5072 = cnt[6] ? _GEN_5062 : _GEN_5052; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5073 = cnt[6] ? _GEN_5063 : _GEN_5053; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_5074 = cnt[6] ? _GEN_5064 : _GEN_5054; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_5075 = cnt[6] ? _GEN_5065 : _GEN_4910; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5076 = _GEN_145 | _GEN_5066; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5077 = _GEN_146 | _GEN_5067; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5078 = _GEN_147 | _GEN_5068; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5079 = _GEN_148 | _GEN_5069; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5080 = 2'h0 == opidx ? 5'hc : _GEN_5070; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5081 = 2'h1 == opidx ? 5'hc : _GEN_5071; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5082 = 2'h2 == opidx ? 5'hc : _GEN_5072; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5083 = 2'h3 == opidx ? 5'hc : _GEN_5073; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_5084 = _T_122 ? _cnt_T : _GEN_5074; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_5085 = _T_122 ? _GEN_1349 : _GEN_4911; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_5086 = cnt[7] ? _GEN_5076 : _GEN_5066; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5087 = cnt[7] ? _GEN_5077 : _GEN_5067; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5088 = cnt[7] ? _GEN_5078 : _GEN_5068; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5089 = cnt[7] ? _GEN_5079 : _GEN_5069; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5090 = cnt[7] ? _GEN_5080 : _GEN_5070; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5091 = cnt[7] ? _GEN_5081 : _GEN_5071; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5092 = cnt[7] ? _GEN_5082 : _GEN_5072; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5093 = cnt[7] ? _GEN_5083 : _GEN_5073; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_5094 = cnt[7] ? _GEN_5084 : _GEN_5074; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_5095 = cnt[7] ? _GEN_5085 : _GEN_4911; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5096 = _GEN_145 | _GEN_5086; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5097 = _GEN_146 | _GEN_5087; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5098 = _GEN_147 | _GEN_5088; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5099 = _GEN_148 | _GEN_5089; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5100 = 2'h0 == opidx ? 5'hd : _GEN_5090; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5101 = 2'h1 == opidx ? 5'hd : _GEN_5091; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5102 = 2'h2 == opidx ? 5'hd : _GEN_5092; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5103 = 2'h3 == opidx ? 5'hd : _GEN_5093; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_5104 = _T_122 ? _cnt_T : _GEN_5094; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_5105 = _T_122 ? _GEN_1349 : _GEN_4912; // @[NulCtrlMP.scala 353:36 355:17]
  wire  _GEN_5106 = cnt[8] ? _GEN_5096 : _GEN_5086; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5107 = cnt[8] ? _GEN_5097 : _GEN_5087; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5108 = cnt[8] ? _GEN_5098 : _GEN_5088; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_5109 = cnt[8] ? _GEN_5099 : _GEN_5089; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5110 = cnt[8] ? _GEN_5100 : _GEN_5090; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5111 = cnt[8] ? _GEN_5101 : _GEN_5091; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5112 = cnt[8] ? _GEN_5102 : _GEN_5092; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_5113 = cnt[8] ? _GEN_5103 : _GEN_5093; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_5114 = cnt[8] ? _GEN_5104 : _GEN_5094; // @[NulCtrlMP.scala 408:32]
  wire [63:0] _GEN_5115 = cnt[8] ? _GEN_5105 : _GEN_4912; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_5116 = io_tx_ready ? _cnt_T : _GEN_5114; // @[NulCtrlMP.scala 827:31 828:21]
  wire  _GEN_5117 = cnt[9] | _GEN_1102; // @[NulCtrlMP.scala 824:22 825:25]
  wire [7:0] _GEN_5118 = cnt[9] ? _io_tx_bits_T : _GEN_1103; // @[NulCtrlMP.scala 824:22 826:24]
  wire [128:0] _GEN_5119 = cnt[9] ? _GEN_5116 : _GEN_5114; // @[NulCtrlMP.scala 824:22]
  wire [11:0] _T_463 = {opoff, 9'h0}; // @[NulCtrlMP.scala 831:61]
  wire [63:0] _GEN_9872 = {{52'd0}, _T_463}; // @[NulCtrlMP.scala 831:52]
  wire [63:0] _T_464 = pg_base_addr2 | _GEN_9872; // @[NulCtrlMP.scala 831:52]
  wire  _GEN_5120 = _GEN_145 | _GEN_4914; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_5121 = _GEN_146 | _GEN_4915; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_5122 = _GEN_147 | _GEN_4916; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_5123 = _GEN_148 | _GEN_4917; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_5124 = 2'h0 == opidx ? 5'h5 : _GEN_5110; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_5125 = 2'h1 == opidx ? 5'h5 : _GEN_5111; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_5126 = 2'h2 == opidx ? 5'h5 : _GEN_5112; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_5127 = 2'h3 == opidx ? 5'h5 : _GEN_5113; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_5128 = 2'h0 == opidx ? _T_464 : _GEN_4918; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_5129 = 2'h1 == opidx ? _T_464 : _GEN_4919; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_5130 = 2'h2 == opidx ? _T_464 : _GEN_4920; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_5131 = 2'h3 == opidx ? _T_464 : _GEN_4921; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_5132 = ~_GEN_1128 ? _cnt_T : _GEN_5119; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_5133 = cnt[10] ? _GEN_5120 : _GEN_4914; // @[NulCtrlMP.scala 831:23]
  wire  _GEN_5134 = cnt[10] ? _GEN_5121 : _GEN_4915; // @[NulCtrlMP.scala 831:23]
  wire  _GEN_5135 = cnt[10] ? _GEN_5122 : _GEN_4916; // @[NulCtrlMP.scala 831:23]
  wire  _GEN_5136 = cnt[10] ? _GEN_5123 : _GEN_4917; // @[NulCtrlMP.scala 831:23]
  wire [4:0] _GEN_5137 = cnt[10] ? _GEN_5124 : _GEN_5110; // @[NulCtrlMP.scala 831:23]
  wire [4:0] _GEN_5138 = cnt[10] ? _GEN_5125 : _GEN_5111; // @[NulCtrlMP.scala 831:23]
  wire [4:0] _GEN_5139 = cnt[10] ? _GEN_5126 : _GEN_5112; // @[NulCtrlMP.scala 831:23]
  wire [4:0] _GEN_5140 = cnt[10] ? _GEN_5127 : _GEN_5113; // @[NulCtrlMP.scala 831:23]
  wire [63:0] _GEN_5141 = cnt[10] ? _GEN_5128 : _GEN_4918; // @[NulCtrlMP.scala 831:23]
  wire [63:0] _GEN_5142 = cnt[10] ? _GEN_5129 : _GEN_4919; // @[NulCtrlMP.scala 831:23]
  wire [63:0] _GEN_5143 = cnt[10] ? _GEN_5130 : _GEN_4920; // @[NulCtrlMP.scala 831:23]
  wire [63:0] _GEN_5144 = cnt[10] ? _GEN_5131 : _GEN_4921; // @[NulCtrlMP.scala 831:23]
  wire [128:0] _GEN_5145 = cnt[10] ? _GEN_5132 : _GEN_5119; // @[NulCtrlMP.scala 831:23]
  wire  _GEN_5146 = _GEN_145 | _GEN_4922; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5147 = _GEN_146 | _GEN_4923; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5148 = _GEN_147 | _GEN_4924; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5149 = _GEN_148 | _GEN_4925; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_5150 = 2'h0 == opidx ? 32'h2b303 : _GEN_4926; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5151 = 2'h1 == opidx ? 32'h2b303 : _GEN_4927; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5152 = 2'h2 == opidx ? 32'h2b303 : _GEN_4928; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5153 = 2'h3 == opidx ? 32'h2b303 : _GEN_4929; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_5154 = _GEN_1180 ? _cnt_T : _GEN_5145; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_5155 = cnt[11] ? _GEN_5146 : _GEN_4922; // @[NulCtrlMP.scala 832:23]
  wire  _GEN_5156 = cnt[11] ? _GEN_5147 : _GEN_4923; // @[NulCtrlMP.scala 832:23]
  wire  _GEN_5157 = cnt[11] ? _GEN_5148 : _GEN_4924; // @[NulCtrlMP.scala 832:23]
  wire  _GEN_5158 = cnt[11] ? _GEN_5149 : _GEN_4925; // @[NulCtrlMP.scala 832:23]
  wire [31:0] _GEN_5159 = cnt[11] ? _GEN_5150 : _GEN_4926; // @[NulCtrlMP.scala 832:23]
  wire [31:0] _GEN_5160 = cnt[11] ? _GEN_5151 : _GEN_4927; // @[NulCtrlMP.scala 832:23]
  wire [31:0] _GEN_5161 = cnt[11] ? _GEN_5152 : _GEN_4928; // @[NulCtrlMP.scala 832:23]
  wire [31:0] _GEN_5162 = cnt[11] ? _GEN_5153 : _GEN_4929; // @[NulCtrlMP.scala 832:23]
  wire [128:0] _GEN_5163 = cnt[11] ? _GEN_5154 : _GEN_5145; // @[NulCtrlMP.scala 832:23]
  wire  _GEN_5164 = _GEN_145 | _GEN_5155; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5165 = _GEN_146 | _GEN_5156; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5166 = _GEN_147 | _GEN_5157; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5167 = _GEN_148 | _GEN_5158; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_5168 = 2'h0 == opidx ? 32'h82b383 : _GEN_5159; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5169 = 2'h1 == opidx ? 32'h82b383 : _GEN_5160; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5170 = 2'h2 == opidx ? 32'h82b383 : _GEN_5161; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5171 = 2'h3 == opidx ? 32'h82b383 : _GEN_5162; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_5172 = _GEN_1180 ? _cnt_T : _GEN_5163; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_5173 = cnt[12] ? _GEN_5164 : _GEN_5155; // @[NulCtrlMP.scala 833:23]
  wire  _GEN_5174 = cnt[12] ? _GEN_5165 : _GEN_5156; // @[NulCtrlMP.scala 833:23]
  wire  _GEN_5175 = cnt[12] ? _GEN_5166 : _GEN_5157; // @[NulCtrlMP.scala 833:23]
  wire  _GEN_5176 = cnt[12] ? _GEN_5167 : _GEN_5158; // @[NulCtrlMP.scala 833:23]
  wire [31:0] _GEN_5177 = cnt[12] ? _GEN_5168 : _GEN_5159; // @[NulCtrlMP.scala 833:23]
  wire [31:0] _GEN_5178 = cnt[12] ? _GEN_5169 : _GEN_5160; // @[NulCtrlMP.scala 833:23]
  wire [31:0] _GEN_5179 = cnt[12] ? _GEN_5170 : _GEN_5161; // @[NulCtrlMP.scala 833:23]
  wire [31:0] _GEN_5180 = cnt[12] ? _GEN_5171 : _GEN_5162; // @[NulCtrlMP.scala 833:23]
  wire [128:0] _GEN_5181 = cnt[12] ? _GEN_5172 : _GEN_5163; // @[NulCtrlMP.scala 833:23]
  wire  _GEN_5182 = _GEN_145 | _GEN_5173; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5183 = _GEN_146 | _GEN_5174; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5184 = _GEN_147 | _GEN_5175; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5185 = _GEN_148 | _GEN_5176; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_5186 = 2'h0 == opidx ? 32'h102b403 : _GEN_5177; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5187 = 2'h1 == opidx ? 32'h102b403 : _GEN_5178; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5188 = 2'h2 == opidx ? 32'h102b403 : _GEN_5179; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5189 = 2'h3 == opidx ? 32'h102b403 : _GEN_5180; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_5190 = _GEN_1180 ? _cnt_T : _GEN_5181; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_5191 = cnt[13] ? _GEN_5182 : _GEN_5173; // @[NulCtrlMP.scala 834:23]
  wire  _GEN_5192 = cnt[13] ? _GEN_5183 : _GEN_5174; // @[NulCtrlMP.scala 834:23]
  wire  _GEN_5193 = cnt[13] ? _GEN_5184 : _GEN_5175; // @[NulCtrlMP.scala 834:23]
  wire  _GEN_5194 = cnt[13] ? _GEN_5185 : _GEN_5176; // @[NulCtrlMP.scala 834:23]
  wire [31:0] _GEN_5195 = cnt[13] ? _GEN_5186 : _GEN_5177; // @[NulCtrlMP.scala 834:23]
  wire [31:0] _GEN_5196 = cnt[13] ? _GEN_5187 : _GEN_5178; // @[NulCtrlMP.scala 834:23]
  wire [31:0] _GEN_5197 = cnt[13] ? _GEN_5188 : _GEN_5179; // @[NulCtrlMP.scala 834:23]
  wire [31:0] _GEN_5198 = cnt[13] ? _GEN_5189 : _GEN_5180; // @[NulCtrlMP.scala 834:23]
  wire [128:0] _GEN_5199 = cnt[13] ? _GEN_5190 : _GEN_5181; // @[NulCtrlMP.scala 834:23]
  wire  _GEN_5200 = _GEN_145 | _GEN_5191; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5201 = _GEN_146 | _GEN_5192; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5202 = _GEN_147 | _GEN_5193; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5203 = _GEN_148 | _GEN_5194; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_5204 = 2'h0 == opidx ? 32'h182b483 : _GEN_5195; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5205 = 2'h1 == opidx ? 32'h182b483 : _GEN_5196; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5206 = 2'h2 == opidx ? 32'h182b483 : _GEN_5197; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5207 = 2'h3 == opidx ? 32'h182b483 : _GEN_5198; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_5208 = _GEN_1180 ? _cnt_T : _GEN_5199; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_5209 = cnt[14] ? _GEN_5200 : _GEN_5191; // @[NulCtrlMP.scala 835:23]
  wire  _GEN_5210 = cnt[14] ? _GEN_5201 : _GEN_5192; // @[NulCtrlMP.scala 835:23]
  wire  _GEN_5211 = cnt[14] ? _GEN_5202 : _GEN_5193; // @[NulCtrlMP.scala 835:23]
  wire  _GEN_5212 = cnt[14] ? _GEN_5203 : _GEN_5194; // @[NulCtrlMP.scala 835:23]
  wire [31:0] _GEN_5213 = cnt[14] ? _GEN_5204 : _GEN_5195; // @[NulCtrlMP.scala 835:23]
  wire [31:0] _GEN_5214 = cnt[14] ? _GEN_5205 : _GEN_5196; // @[NulCtrlMP.scala 835:23]
  wire [31:0] _GEN_5215 = cnt[14] ? _GEN_5206 : _GEN_5197; // @[NulCtrlMP.scala 835:23]
  wire [31:0] _GEN_5216 = cnt[14] ? _GEN_5207 : _GEN_5198; // @[NulCtrlMP.scala 835:23]
  wire [128:0] _GEN_5217 = cnt[14] ? _GEN_5208 : _GEN_5199; // @[NulCtrlMP.scala 835:23]
  wire  _GEN_5218 = _GEN_145 | _GEN_5209; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5219 = _GEN_146 | _GEN_5210; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5220 = _GEN_147 | _GEN_5211; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5221 = _GEN_148 | _GEN_5212; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_5222 = 2'h0 == opidx ? 32'h202b503 : _GEN_5213; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5223 = 2'h1 == opidx ? 32'h202b503 : _GEN_5214; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5224 = 2'h2 == opidx ? 32'h202b503 : _GEN_5215; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5225 = 2'h3 == opidx ? 32'h202b503 : _GEN_5216; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_5226 = _GEN_1180 ? _cnt_T : _GEN_5217; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_5227 = cnt[15] ? _GEN_5218 : _GEN_5209; // @[NulCtrlMP.scala 836:23]
  wire  _GEN_5228 = cnt[15] ? _GEN_5219 : _GEN_5210; // @[NulCtrlMP.scala 836:23]
  wire  _GEN_5229 = cnt[15] ? _GEN_5220 : _GEN_5211; // @[NulCtrlMP.scala 836:23]
  wire  _GEN_5230 = cnt[15] ? _GEN_5221 : _GEN_5212; // @[NulCtrlMP.scala 836:23]
  wire [31:0] _GEN_5231 = cnt[15] ? _GEN_5222 : _GEN_5213; // @[NulCtrlMP.scala 836:23]
  wire [31:0] _GEN_5232 = cnt[15] ? _GEN_5223 : _GEN_5214; // @[NulCtrlMP.scala 836:23]
  wire [31:0] _GEN_5233 = cnt[15] ? _GEN_5224 : _GEN_5215; // @[NulCtrlMP.scala 836:23]
  wire [31:0] _GEN_5234 = cnt[15] ? _GEN_5225 : _GEN_5216; // @[NulCtrlMP.scala 836:23]
  wire [128:0] _GEN_5235 = cnt[15] ? _GEN_5226 : _GEN_5217; // @[NulCtrlMP.scala 836:23]
  wire  _GEN_5236 = _GEN_145 | _GEN_5227; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5237 = _GEN_146 | _GEN_5228; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5238 = _GEN_147 | _GEN_5229; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5239 = _GEN_148 | _GEN_5230; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_5240 = 2'h0 == opidx ? 32'h282b583 : _GEN_5231; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5241 = 2'h1 == opidx ? 32'h282b583 : _GEN_5232; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5242 = 2'h2 == opidx ? 32'h282b583 : _GEN_5233; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5243 = 2'h3 == opidx ? 32'h282b583 : _GEN_5234; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_5244 = _GEN_1180 ? _cnt_T : _GEN_5235; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_5245 = cnt[16] ? _GEN_5236 : _GEN_5227; // @[NulCtrlMP.scala 837:23]
  wire  _GEN_5246 = cnt[16] ? _GEN_5237 : _GEN_5228; // @[NulCtrlMP.scala 837:23]
  wire  _GEN_5247 = cnt[16] ? _GEN_5238 : _GEN_5229; // @[NulCtrlMP.scala 837:23]
  wire  _GEN_5248 = cnt[16] ? _GEN_5239 : _GEN_5230; // @[NulCtrlMP.scala 837:23]
  wire [31:0] _GEN_5249 = cnt[16] ? _GEN_5240 : _GEN_5231; // @[NulCtrlMP.scala 837:23]
  wire [31:0] _GEN_5250 = cnt[16] ? _GEN_5241 : _GEN_5232; // @[NulCtrlMP.scala 837:23]
  wire [31:0] _GEN_5251 = cnt[16] ? _GEN_5242 : _GEN_5233; // @[NulCtrlMP.scala 837:23]
  wire [31:0] _GEN_5252 = cnt[16] ? _GEN_5243 : _GEN_5234; // @[NulCtrlMP.scala 837:23]
  wire [128:0] _GEN_5253 = cnt[16] ? _GEN_5244 : _GEN_5235; // @[NulCtrlMP.scala 837:23]
  wire  _GEN_5254 = _GEN_145 | _GEN_5245; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5255 = _GEN_146 | _GEN_5246; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5256 = _GEN_147 | _GEN_5247; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5257 = _GEN_148 | _GEN_5248; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_5258 = 2'h0 == opidx ? 32'h302b603 : _GEN_5249; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5259 = 2'h1 == opidx ? 32'h302b603 : _GEN_5250; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5260 = 2'h2 == opidx ? 32'h302b603 : _GEN_5251; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5261 = 2'h3 == opidx ? 32'h302b603 : _GEN_5252; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_5262 = _GEN_1180 ? _cnt_T : _GEN_5253; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_5263 = cnt[17] ? _GEN_5254 : _GEN_5245; // @[NulCtrlMP.scala 838:23]
  wire  _GEN_5264 = cnt[17] ? _GEN_5255 : _GEN_5246; // @[NulCtrlMP.scala 838:23]
  wire  _GEN_5265 = cnt[17] ? _GEN_5256 : _GEN_5247; // @[NulCtrlMP.scala 838:23]
  wire  _GEN_5266 = cnt[17] ? _GEN_5257 : _GEN_5248; // @[NulCtrlMP.scala 838:23]
  wire [31:0] _GEN_5267 = cnt[17] ? _GEN_5258 : _GEN_5249; // @[NulCtrlMP.scala 838:23]
  wire [31:0] _GEN_5268 = cnt[17] ? _GEN_5259 : _GEN_5250; // @[NulCtrlMP.scala 838:23]
  wire [31:0] _GEN_5269 = cnt[17] ? _GEN_5260 : _GEN_5251; // @[NulCtrlMP.scala 838:23]
  wire [31:0] _GEN_5270 = cnt[17] ? _GEN_5261 : _GEN_5252; // @[NulCtrlMP.scala 838:23]
  wire [128:0] _GEN_5271 = cnt[17] ? _GEN_5262 : _GEN_5253; // @[NulCtrlMP.scala 838:23]
  wire  _GEN_5272 = _GEN_145 | _GEN_5263; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5273 = _GEN_146 | _GEN_5264; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5274 = _GEN_147 | _GEN_5265; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5275 = _GEN_148 | _GEN_5266; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_5276 = 2'h0 == opidx ? 32'h382b683 : _GEN_5267; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5277 = 2'h1 == opidx ? 32'h382b683 : _GEN_5268; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5278 = 2'h2 == opidx ? 32'h382b683 : _GEN_5269; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5279 = 2'h3 == opidx ? 32'h382b683 : _GEN_5270; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_5280 = _GEN_1180 ? _cnt_T : _GEN_5271; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_5281 = cnt[18] ? _GEN_5272 : _GEN_5263; // @[NulCtrlMP.scala 839:23]
  wire  _GEN_5282 = cnt[18] ? _GEN_5273 : _GEN_5264; // @[NulCtrlMP.scala 839:23]
  wire  _GEN_5283 = cnt[18] ? _GEN_5274 : _GEN_5265; // @[NulCtrlMP.scala 839:23]
  wire  _GEN_5284 = cnt[18] ? _GEN_5275 : _GEN_5266; // @[NulCtrlMP.scala 839:23]
  wire [31:0] _GEN_5285 = cnt[18] ? _GEN_5276 : _GEN_5267; // @[NulCtrlMP.scala 839:23]
  wire [31:0] _GEN_5286 = cnt[18] ? _GEN_5277 : _GEN_5268; // @[NulCtrlMP.scala 839:23]
  wire [31:0] _GEN_5287 = cnt[18] ? _GEN_5278 : _GEN_5269; // @[NulCtrlMP.scala 839:23]
  wire [31:0] _GEN_5288 = cnt[18] ? _GEN_5279 : _GEN_5270; // @[NulCtrlMP.scala 839:23]
  wire [128:0] _GEN_5289 = cnt[18] ? _GEN_5280 : _GEN_5271; // @[NulCtrlMP.scala 839:23]
  wire  _GEN_5290 = _GEN_145 | _GEN_5281; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5291 = _GEN_146 | _GEN_5282; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5292 = _GEN_147 | _GEN_5283; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_5293 = _GEN_148 | _GEN_5284; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_5294 = 2'h0 == opidx ? 32'h4028293 : _GEN_5285; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5295 = 2'h1 == opidx ? 32'h4028293 : _GEN_5286; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5296 = 2'h2 == opidx ? 32'h4028293 : _GEN_5287; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_5297 = 2'h3 == opidx ? 32'h4028293 : _GEN_5288; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_5298 = _GEN_1180 ? _cnt_T : _GEN_5289; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_5299 = cnt[19] ? _GEN_5290 : _GEN_5281; // @[NulCtrlMP.scala 840:23]
  wire  _GEN_5300 = cnt[19] ? _GEN_5291 : _GEN_5282; // @[NulCtrlMP.scala 840:23]
  wire  _GEN_5301 = cnt[19] ? _GEN_5292 : _GEN_5283; // @[NulCtrlMP.scala 840:23]
  wire  _GEN_5302 = cnt[19] ? _GEN_5293 : _GEN_5284; // @[NulCtrlMP.scala 840:23]
  wire [31:0] _GEN_5303 = cnt[19] ? _GEN_5294 : _GEN_5285; // @[NulCtrlMP.scala 840:23]
  wire [31:0] _GEN_5304 = cnt[19] ? _GEN_5295 : _GEN_5286; // @[NulCtrlMP.scala 840:23]
  wire [31:0] _GEN_5305 = cnt[19] ? _GEN_5296 : _GEN_5287; // @[NulCtrlMP.scala 840:23]
  wire [31:0] _GEN_5306 = cnt[19] ? _GEN_5297 : _GEN_5288; // @[NulCtrlMP.scala 840:23]
  wire [128:0] _GEN_5307 = cnt[19] ? _GEN_5298 : _GEN_5289; // @[NulCtrlMP.scala 840:23]
  wire  _GEN_5308 = _GEN_145 | _GEN_4930; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_5309 = _GEN_146 | _GEN_4931; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_5310 = _GEN_147 | _GEN_4932; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_5311 = _GEN_148 | _GEN_4933; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_5312 = ~_GEN_1252 ? _cnt_T : _GEN_5307; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_5313 = cnt[20] ? _GEN_5308 : _GEN_4930; // @[NulCtrlMP.scala 841:23]
  wire  _GEN_5314 = cnt[20] ? _GEN_5309 : _GEN_4931; // @[NulCtrlMP.scala 841:23]
  wire  _GEN_5315 = cnt[20] ? _GEN_5310 : _GEN_4932; // @[NulCtrlMP.scala 841:23]
  wire  _GEN_5316 = cnt[20] ? _GEN_5311 : _GEN_4933; // @[NulCtrlMP.scala 841:23]
  wire [128:0] _GEN_5317 = cnt[20] ? _GEN_5312 : _GEN_5307; // @[NulCtrlMP.scala 841:23]
  wire [9:0] _T_479 = {{1'd0}, pgbuf_cpu_pos[11:3]}; // @[NulCtrlMP.scala 843:77]
  wire  _GEN_5318 = _GEN_145 | _GEN_5106; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5319 = _GEN_146 | _GEN_5107; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5320 = _GEN_147 | _GEN_5108; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5321 = _GEN_148 | _GEN_5109; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5322 = 2'h0 == opidx ? 5'h6 : _GEN_5137; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5323 = 2'h1 == opidx ? 5'h6 : _GEN_5138; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5324 = 2'h2 == opidx ? 5'h6 : _GEN_5139; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5325 = 2'h3 == opidx ? 5'h6 : _GEN_5140; // @[NulCtrlMP.scala 352:{28,28}]
  wire [63:0] _GEN_5326 = 6'h0 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_0; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5327 = 6'h1 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_1; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5328 = 6'h2 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_2; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5329 = 6'h3 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_3; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5330 = 6'h4 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_4; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5331 = 6'h5 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_5; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5332 = 6'h6 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_6; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5333 = 6'h7 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_7; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5334 = 6'h8 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_8; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5335 = 6'h9 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_9; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5336 = 6'ha == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_10; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5337 = 6'hb == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_11; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5338 = 6'hc == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_12; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5339 = 6'hd == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_13; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5340 = 6'he == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_14; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5341 = 6'hf == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_15; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5342 = 6'h10 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_16; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5343 = 6'h11 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_17; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5344 = 6'h12 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_18; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5345 = 6'h13 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_19; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5346 = 6'h14 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_20; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5347 = 6'h15 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_21; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5348 = 6'h16 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_22; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5349 = 6'h17 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_23; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5350 = 6'h18 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_24; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5351 = 6'h19 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_25; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5352 = 6'h1a == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_26; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5353 = 6'h1b == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_27; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5354 = 6'h1c == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_28; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5355 = 6'h1d == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_29; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5356 = 6'h1e == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_30; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5357 = 6'h1f == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_31; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5358 = 6'h20 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_32; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5359 = 6'h21 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_33; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5360 = 6'h22 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_34; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5361 = 6'h23 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_35; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5362 = 6'h24 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_36; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5363 = 6'h25 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_37; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5364 = 6'h26 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_38; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5365 = 6'h27 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_39; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5366 = 6'h28 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_40; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5367 = 6'h29 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_41; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5368 = 6'h2a == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_42; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5369 = 6'h2b == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_43; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5370 = 6'h2c == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_44; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5371 = 6'h2d == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_45; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5372 = 6'h2e == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_46; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5373 = 6'h2f == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_47; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5374 = 6'h30 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_48; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5375 = 6'h31 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_49; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5376 = 6'h32 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_50; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5377 = 6'h33 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_51; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5378 = 6'h34 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_52; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5379 = 6'h35 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_53; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5380 = 6'h36 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_54; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5381 = 6'h37 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_55; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5382 = 6'h38 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_56; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5383 = 6'h39 == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_57; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5384 = 6'h3a == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_58; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5385 = 6'h3b == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_59; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5386 = 6'h3c == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_60; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5387 = 6'h3d == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_61; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5388 = 6'h3e == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_62; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [63:0] _GEN_5389 = 6'h3f == _T_479[5:0] ? _GEN_1349 : pgbuf_div8_63; // @[NulCtrlMP.scala 355:{17,17} 818:29]
  wire [128:0] _GEN_5390 = _T_122 ? _cnt_T : _GEN_5317; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_5391 = _T_122 ? _GEN_5326 : pgbuf_div8_0; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5392 = _T_122 ? _GEN_5327 : pgbuf_div8_1; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5393 = _T_122 ? _GEN_5328 : pgbuf_div8_2; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5394 = _T_122 ? _GEN_5329 : pgbuf_div8_3; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5395 = _T_122 ? _GEN_5330 : pgbuf_div8_4; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5396 = _T_122 ? _GEN_5331 : pgbuf_div8_5; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5397 = _T_122 ? _GEN_5332 : pgbuf_div8_6; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5398 = _T_122 ? _GEN_5333 : pgbuf_div8_7; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5399 = _T_122 ? _GEN_5334 : pgbuf_div8_8; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5400 = _T_122 ? _GEN_5335 : pgbuf_div8_9; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5401 = _T_122 ? _GEN_5336 : pgbuf_div8_10; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5402 = _T_122 ? _GEN_5337 : pgbuf_div8_11; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5403 = _T_122 ? _GEN_5338 : pgbuf_div8_12; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5404 = _T_122 ? _GEN_5339 : pgbuf_div8_13; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5405 = _T_122 ? _GEN_5340 : pgbuf_div8_14; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5406 = _T_122 ? _GEN_5341 : pgbuf_div8_15; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5407 = _T_122 ? _GEN_5342 : pgbuf_div8_16; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5408 = _T_122 ? _GEN_5343 : pgbuf_div8_17; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5409 = _T_122 ? _GEN_5344 : pgbuf_div8_18; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5410 = _T_122 ? _GEN_5345 : pgbuf_div8_19; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5411 = _T_122 ? _GEN_5346 : pgbuf_div8_20; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5412 = _T_122 ? _GEN_5347 : pgbuf_div8_21; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5413 = _T_122 ? _GEN_5348 : pgbuf_div8_22; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5414 = _T_122 ? _GEN_5349 : pgbuf_div8_23; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5415 = _T_122 ? _GEN_5350 : pgbuf_div8_24; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5416 = _T_122 ? _GEN_5351 : pgbuf_div8_25; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5417 = _T_122 ? _GEN_5352 : pgbuf_div8_26; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5418 = _T_122 ? _GEN_5353 : pgbuf_div8_27; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5419 = _T_122 ? _GEN_5354 : pgbuf_div8_28; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5420 = _T_122 ? _GEN_5355 : pgbuf_div8_29; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5421 = _T_122 ? _GEN_5356 : pgbuf_div8_30; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5422 = _T_122 ? _GEN_5357 : pgbuf_div8_31; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5423 = _T_122 ? _GEN_5358 : pgbuf_div8_32; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5424 = _T_122 ? _GEN_5359 : pgbuf_div8_33; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5425 = _T_122 ? _GEN_5360 : pgbuf_div8_34; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5426 = _T_122 ? _GEN_5361 : pgbuf_div8_35; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5427 = _T_122 ? _GEN_5362 : pgbuf_div8_36; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5428 = _T_122 ? _GEN_5363 : pgbuf_div8_37; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5429 = _T_122 ? _GEN_5364 : pgbuf_div8_38; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5430 = _T_122 ? _GEN_5365 : pgbuf_div8_39; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5431 = _T_122 ? _GEN_5366 : pgbuf_div8_40; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5432 = _T_122 ? _GEN_5367 : pgbuf_div8_41; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5433 = _T_122 ? _GEN_5368 : pgbuf_div8_42; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5434 = _T_122 ? _GEN_5369 : pgbuf_div8_43; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5435 = _T_122 ? _GEN_5370 : pgbuf_div8_44; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5436 = _T_122 ? _GEN_5371 : pgbuf_div8_45; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5437 = _T_122 ? _GEN_5372 : pgbuf_div8_46; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5438 = _T_122 ? _GEN_5373 : pgbuf_div8_47; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5439 = _T_122 ? _GEN_5374 : pgbuf_div8_48; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5440 = _T_122 ? _GEN_5375 : pgbuf_div8_49; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5441 = _T_122 ? _GEN_5376 : pgbuf_div8_50; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5442 = _T_122 ? _GEN_5377 : pgbuf_div8_51; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5443 = _T_122 ? _GEN_5378 : pgbuf_div8_52; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5444 = _T_122 ? _GEN_5379 : pgbuf_div8_53; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5445 = _T_122 ? _GEN_5380 : pgbuf_div8_54; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5446 = _T_122 ? _GEN_5381 : pgbuf_div8_55; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5447 = _T_122 ? _GEN_5382 : pgbuf_div8_56; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5448 = _T_122 ? _GEN_5383 : pgbuf_div8_57; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5449 = _T_122 ? _GEN_5384 : pgbuf_div8_58; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5450 = _T_122 ? _GEN_5385 : pgbuf_div8_59; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5451 = _T_122 ? _GEN_5386 : pgbuf_div8_60; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5452 = _T_122 ? _GEN_5387 : pgbuf_div8_61; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5453 = _T_122 ? _GEN_5388 : pgbuf_div8_62; // @[NulCtrlMP.scala 353:36 818:29]
  wire [63:0] _GEN_5454 = _T_122 ? _GEN_5389 : pgbuf_div8_63; // @[NulCtrlMP.scala 353:36 818:29]
  wire  _GEN_5455 = cnt[21] ? _GEN_5318 : _GEN_5106; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_5456 = cnt[21] ? _GEN_5319 : _GEN_5107; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_5457 = cnt[21] ? _GEN_5320 : _GEN_5108; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_5458 = cnt[21] ? _GEN_5321 : _GEN_5109; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5459 = cnt[21] ? _GEN_5322 : _GEN_5137; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5460 = cnt[21] ? _GEN_5323 : _GEN_5138; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5461 = cnt[21] ? _GEN_5324 : _GEN_5139; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5462 = cnt[21] ? _GEN_5325 : _GEN_5140; // @[NulCtrlMP.scala 843:29]
  wire [128:0] _GEN_5463 = cnt[21] ? _GEN_5390 : _GEN_5317; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5464 = cnt[21] ? _GEN_5391 : pgbuf_div8_0; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5465 = cnt[21] ? _GEN_5392 : pgbuf_div8_1; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5466 = cnt[21] ? _GEN_5393 : pgbuf_div8_2; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5467 = cnt[21] ? _GEN_5394 : pgbuf_div8_3; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5468 = cnt[21] ? _GEN_5395 : pgbuf_div8_4; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5469 = cnt[21] ? _GEN_5396 : pgbuf_div8_5; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5470 = cnt[21] ? _GEN_5397 : pgbuf_div8_6; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5471 = cnt[21] ? _GEN_5398 : pgbuf_div8_7; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5472 = cnt[21] ? _GEN_5399 : pgbuf_div8_8; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5473 = cnt[21] ? _GEN_5400 : pgbuf_div8_9; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5474 = cnt[21] ? _GEN_5401 : pgbuf_div8_10; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5475 = cnt[21] ? _GEN_5402 : pgbuf_div8_11; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5476 = cnt[21] ? _GEN_5403 : pgbuf_div8_12; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5477 = cnt[21] ? _GEN_5404 : pgbuf_div8_13; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5478 = cnt[21] ? _GEN_5405 : pgbuf_div8_14; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5479 = cnt[21] ? _GEN_5406 : pgbuf_div8_15; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5480 = cnt[21] ? _GEN_5407 : pgbuf_div8_16; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5481 = cnt[21] ? _GEN_5408 : pgbuf_div8_17; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5482 = cnt[21] ? _GEN_5409 : pgbuf_div8_18; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5483 = cnt[21] ? _GEN_5410 : pgbuf_div8_19; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5484 = cnt[21] ? _GEN_5411 : pgbuf_div8_20; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5485 = cnt[21] ? _GEN_5412 : pgbuf_div8_21; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5486 = cnt[21] ? _GEN_5413 : pgbuf_div8_22; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5487 = cnt[21] ? _GEN_5414 : pgbuf_div8_23; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5488 = cnt[21] ? _GEN_5415 : pgbuf_div8_24; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5489 = cnt[21] ? _GEN_5416 : pgbuf_div8_25; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5490 = cnt[21] ? _GEN_5417 : pgbuf_div8_26; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5491 = cnt[21] ? _GEN_5418 : pgbuf_div8_27; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5492 = cnt[21] ? _GEN_5419 : pgbuf_div8_28; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5493 = cnt[21] ? _GEN_5420 : pgbuf_div8_29; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5494 = cnt[21] ? _GEN_5421 : pgbuf_div8_30; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5495 = cnt[21] ? _GEN_5422 : pgbuf_div8_31; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5496 = cnt[21] ? _GEN_5423 : pgbuf_div8_32; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5497 = cnt[21] ? _GEN_5424 : pgbuf_div8_33; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5498 = cnt[21] ? _GEN_5425 : pgbuf_div8_34; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5499 = cnt[21] ? _GEN_5426 : pgbuf_div8_35; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5500 = cnt[21] ? _GEN_5427 : pgbuf_div8_36; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5501 = cnt[21] ? _GEN_5428 : pgbuf_div8_37; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5502 = cnt[21] ? _GEN_5429 : pgbuf_div8_38; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5503 = cnt[21] ? _GEN_5430 : pgbuf_div8_39; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5504 = cnt[21] ? _GEN_5431 : pgbuf_div8_40; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5505 = cnt[21] ? _GEN_5432 : pgbuf_div8_41; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5506 = cnt[21] ? _GEN_5433 : pgbuf_div8_42; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5507 = cnt[21] ? _GEN_5434 : pgbuf_div8_43; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5508 = cnt[21] ? _GEN_5435 : pgbuf_div8_44; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5509 = cnt[21] ? _GEN_5436 : pgbuf_div8_45; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5510 = cnt[21] ? _GEN_5437 : pgbuf_div8_46; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5511 = cnt[21] ? _GEN_5438 : pgbuf_div8_47; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5512 = cnt[21] ? _GEN_5439 : pgbuf_div8_48; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5513 = cnt[21] ? _GEN_5440 : pgbuf_div8_49; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5514 = cnt[21] ? _GEN_5441 : pgbuf_div8_50; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5515 = cnt[21] ? _GEN_5442 : pgbuf_div8_51; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5516 = cnt[21] ? _GEN_5443 : pgbuf_div8_52; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5517 = cnt[21] ? _GEN_5444 : pgbuf_div8_53; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5518 = cnt[21] ? _GEN_5445 : pgbuf_div8_54; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5519 = cnt[21] ? _GEN_5446 : pgbuf_div8_55; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5520 = cnt[21] ? _GEN_5447 : pgbuf_div8_56; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5521 = cnt[21] ? _GEN_5448 : pgbuf_div8_57; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5522 = cnt[21] ? _GEN_5449 : pgbuf_div8_58; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5523 = cnt[21] ? _GEN_5450 : pgbuf_div8_59; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5524 = cnt[21] ? _GEN_5451 : pgbuf_div8_60; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5525 = cnt[21] ? _GEN_5452 : pgbuf_div8_61; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5526 = cnt[21] ? _GEN_5453 : pgbuf_div8_62; // @[NulCtrlMP.scala 818:29 843:29]
  wire [63:0] _GEN_5527 = cnt[21] ? _GEN_5454 : pgbuf_div8_63; // @[NulCtrlMP.scala 818:29 843:29]
  wire [8:0] _T_486 = pgbuf_cpu_pos[11:3] + 9'h1; // @[NulCtrlMP.scala 843:77]
  wire  _GEN_5528 = _GEN_145 | _GEN_5455; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5529 = _GEN_146 | _GEN_5456; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5530 = _GEN_147 | _GEN_5457; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5531 = _GEN_148 | _GEN_5458; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5532 = 2'h0 == opidx ? 5'h7 : _GEN_5459; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5533 = 2'h1 == opidx ? 5'h7 : _GEN_5460; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5534 = 2'h2 == opidx ? 5'h7 : _GEN_5461; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5535 = 2'h3 == opidx ? 5'h7 : _GEN_5462; // @[NulCtrlMP.scala 352:{28,28}]
  wire [63:0] _GEN_5536 = 6'h0 == _T_486[5:0] ? _GEN_1349 : _GEN_5464; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5537 = 6'h1 == _T_486[5:0] ? _GEN_1349 : _GEN_5465; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5538 = 6'h2 == _T_486[5:0] ? _GEN_1349 : _GEN_5466; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5539 = 6'h3 == _T_486[5:0] ? _GEN_1349 : _GEN_5467; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5540 = 6'h4 == _T_486[5:0] ? _GEN_1349 : _GEN_5468; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5541 = 6'h5 == _T_486[5:0] ? _GEN_1349 : _GEN_5469; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5542 = 6'h6 == _T_486[5:0] ? _GEN_1349 : _GEN_5470; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5543 = 6'h7 == _T_486[5:0] ? _GEN_1349 : _GEN_5471; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5544 = 6'h8 == _T_486[5:0] ? _GEN_1349 : _GEN_5472; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5545 = 6'h9 == _T_486[5:0] ? _GEN_1349 : _GEN_5473; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5546 = 6'ha == _T_486[5:0] ? _GEN_1349 : _GEN_5474; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5547 = 6'hb == _T_486[5:0] ? _GEN_1349 : _GEN_5475; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5548 = 6'hc == _T_486[5:0] ? _GEN_1349 : _GEN_5476; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5549 = 6'hd == _T_486[5:0] ? _GEN_1349 : _GEN_5477; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5550 = 6'he == _T_486[5:0] ? _GEN_1349 : _GEN_5478; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5551 = 6'hf == _T_486[5:0] ? _GEN_1349 : _GEN_5479; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5552 = 6'h10 == _T_486[5:0] ? _GEN_1349 : _GEN_5480; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5553 = 6'h11 == _T_486[5:0] ? _GEN_1349 : _GEN_5481; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5554 = 6'h12 == _T_486[5:0] ? _GEN_1349 : _GEN_5482; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5555 = 6'h13 == _T_486[5:0] ? _GEN_1349 : _GEN_5483; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5556 = 6'h14 == _T_486[5:0] ? _GEN_1349 : _GEN_5484; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5557 = 6'h15 == _T_486[5:0] ? _GEN_1349 : _GEN_5485; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5558 = 6'h16 == _T_486[5:0] ? _GEN_1349 : _GEN_5486; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5559 = 6'h17 == _T_486[5:0] ? _GEN_1349 : _GEN_5487; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5560 = 6'h18 == _T_486[5:0] ? _GEN_1349 : _GEN_5488; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5561 = 6'h19 == _T_486[5:0] ? _GEN_1349 : _GEN_5489; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5562 = 6'h1a == _T_486[5:0] ? _GEN_1349 : _GEN_5490; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5563 = 6'h1b == _T_486[5:0] ? _GEN_1349 : _GEN_5491; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5564 = 6'h1c == _T_486[5:0] ? _GEN_1349 : _GEN_5492; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5565 = 6'h1d == _T_486[5:0] ? _GEN_1349 : _GEN_5493; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5566 = 6'h1e == _T_486[5:0] ? _GEN_1349 : _GEN_5494; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5567 = 6'h1f == _T_486[5:0] ? _GEN_1349 : _GEN_5495; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5568 = 6'h20 == _T_486[5:0] ? _GEN_1349 : _GEN_5496; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5569 = 6'h21 == _T_486[5:0] ? _GEN_1349 : _GEN_5497; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5570 = 6'h22 == _T_486[5:0] ? _GEN_1349 : _GEN_5498; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5571 = 6'h23 == _T_486[5:0] ? _GEN_1349 : _GEN_5499; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5572 = 6'h24 == _T_486[5:0] ? _GEN_1349 : _GEN_5500; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5573 = 6'h25 == _T_486[5:0] ? _GEN_1349 : _GEN_5501; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5574 = 6'h26 == _T_486[5:0] ? _GEN_1349 : _GEN_5502; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5575 = 6'h27 == _T_486[5:0] ? _GEN_1349 : _GEN_5503; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5576 = 6'h28 == _T_486[5:0] ? _GEN_1349 : _GEN_5504; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5577 = 6'h29 == _T_486[5:0] ? _GEN_1349 : _GEN_5505; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5578 = 6'h2a == _T_486[5:0] ? _GEN_1349 : _GEN_5506; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5579 = 6'h2b == _T_486[5:0] ? _GEN_1349 : _GEN_5507; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5580 = 6'h2c == _T_486[5:0] ? _GEN_1349 : _GEN_5508; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5581 = 6'h2d == _T_486[5:0] ? _GEN_1349 : _GEN_5509; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5582 = 6'h2e == _T_486[5:0] ? _GEN_1349 : _GEN_5510; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5583 = 6'h2f == _T_486[5:0] ? _GEN_1349 : _GEN_5511; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5584 = 6'h30 == _T_486[5:0] ? _GEN_1349 : _GEN_5512; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5585 = 6'h31 == _T_486[5:0] ? _GEN_1349 : _GEN_5513; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5586 = 6'h32 == _T_486[5:0] ? _GEN_1349 : _GEN_5514; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5587 = 6'h33 == _T_486[5:0] ? _GEN_1349 : _GEN_5515; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5588 = 6'h34 == _T_486[5:0] ? _GEN_1349 : _GEN_5516; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5589 = 6'h35 == _T_486[5:0] ? _GEN_1349 : _GEN_5517; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5590 = 6'h36 == _T_486[5:0] ? _GEN_1349 : _GEN_5518; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5591 = 6'h37 == _T_486[5:0] ? _GEN_1349 : _GEN_5519; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5592 = 6'h38 == _T_486[5:0] ? _GEN_1349 : _GEN_5520; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5593 = 6'h39 == _T_486[5:0] ? _GEN_1349 : _GEN_5521; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5594 = 6'h3a == _T_486[5:0] ? _GEN_1349 : _GEN_5522; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5595 = 6'h3b == _T_486[5:0] ? _GEN_1349 : _GEN_5523; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5596 = 6'h3c == _T_486[5:0] ? _GEN_1349 : _GEN_5524; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5597 = 6'h3d == _T_486[5:0] ? _GEN_1349 : _GEN_5525; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5598 = 6'h3e == _T_486[5:0] ? _GEN_1349 : _GEN_5526; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5599 = 6'h3f == _T_486[5:0] ? _GEN_1349 : _GEN_5527; // @[NulCtrlMP.scala 355:{17,17}]
  wire [128:0] _GEN_5600 = _T_122 ? _cnt_T : _GEN_5463; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_5601 = _T_122 ? _GEN_5536 : _GEN_5464; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5602 = _T_122 ? _GEN_5537 : _GEN_5465; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5603 = _T_122 ? _GEN_5538 : _GEN_5466; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5604 = _T_122 ? _GEN_5539 : _GEN_5467; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5605 = _T_122 ? _GEN_5540 : _GEN_5468; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5606 = _T_122 ? _GEN_5541 : _GEN_5469; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5607 = _T_122 ? _GEN_5542 : _GEN_5470; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5608 = _T_122 ? _GEN_5543 : _GEN_5471; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5609 = _T_122 ? _GEN_5544 : _GEN_5472; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5610 = _T_122 ? _GEN_5545 : _GEN_5473; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5611 = _T_122 ? _GEN_5546 : _GEN_5474; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5612 = _T_122 ? _GEN_5547 : _GEN_5475; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5613 = _T_122 ? _GEN_5548 : _GEN_5476; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5614 = _T_122 ? _GEN_5549 : _GEN_5477; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5615 = _T_122 ? _GEN_5550 : _GEN_5478; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5616 = _T_122 ? _GEN_5551 : _GEN_5479; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5617 = _T_122 ? _GEN_5552 : _GEN_5480; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5618 = _T_122 ? _GEN_5553 : _GEN_5481; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5619 = _T_122 ? _GEN_5554 : _GEN_5482; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5620 = _T_122 ? _GEN_5555 : _GEN_5483; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5621 = _T_122 ? _GEN_5556 : _GEN_5484; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5622 = _T_122 ? _GEN_5557 : _GEN_5485; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5623 = _T_122 ? _GEN_5558 : _GEN_5486; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5624 = _T_122 ? _GEN_5559 : _GEN_5487; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5625 = _T_122 ? _GEN_5560 : _GEN_5488; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5626 = _T_122 ? _GEN_5561 : _GEN_5489; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5627 = _T_122 ? _GEN_5562 : _GEN_5490; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5628 = _T_122 ? _GEN_5563 : _GEN_5491; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5629 = _T_122 ? _GEN_5564 : _GEN_5492; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5630 = _T_122 ? _GEN_5565 : _GEN_5493; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5631 = _T_122 ? _GEN_5566 : _GEN_5494; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5632 = _T_122 ? _GEN_5567 : _GEN_5495; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5633 = _T_122 ? _GEN_5568 : _GEN_5496; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5634 = _T_122 ? _GEN_5569 : _GEN_5497; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5635 = _T_122 ? _GEN_5570 : _GEN_5498; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5636 = _T_122 ? _GEN_5571 : _GEN_5499; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5637 = _T_122 ? _GEN_5572 : _GEN_5500; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5638 = _T_122 ? _GEN_5573 : _GEN_5501; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5639 = _T_122 ? _GEN_5574 : _GEN_5502; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5640 = _T_122 ? _GEN_5575 : _GEN_5503; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5641 = _T_122 ? _GEN_5576 : _GEN_5504; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5642 = _T_122 ? _GEN_5577 : _GEN_5505; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5643 = _T_122 ? _GEN_5578 : _GEN_5506; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5644 = _T_122 ? _GEN_5579 : _GEN_5507; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5645 = _T_122 ? _GEN_5580 : _GEN_5508; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5646 = _T_122 ? _GEN_5581 : _GEN_5509; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5647 = _T_122 ? _GEN_5582 : _GEN_5510; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5648 = _T_122 ? _GEN_5583 : _GEN_5511; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5649 = _T_122 ? _GEN_5584 : _GEN_5512; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5650 = _T_122 ? _GEN_5585 : _GEN_5513; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5651 = _T_122 ? _GEN_5586 : _GEN_5514; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5652 = _T_122 ? _GEN_5587 : _GEN_5515; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5653 = _T_122 ? _GEN_5588 : _GEN_5516; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5654 = _T_122 ? _GEN_5589 : _GEN_5517; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5655 = _T_122 ? _GEN_5590 : _GEN_5518; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5656 = _T_122 ? _GEN_5591 : _GEN_5519; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5657 = _T_122 ? _GEN_5592 : _GEN_5520; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5658 = _T_122 ? _GEN_5593 : _GEN_5521; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5659 = _T_122 ? _GEN_5594 : _GEN_5522; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5660 = _T_122 ? _GEN_5595 : _GEN_5523; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5661 = _T_122 ? _GEN_5596 : _GEN_5524; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5662 = _T_122 ? _GEN_5597 : _GEN_5525; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5663 = _T_122 ? _GEN_5598 : _GEN_5526; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5664 = _T_122 ? _GEN_5599 : _GEN_5527; // @[NulCtrlMP.scala 353:36]
  wire  _GEN_5665 = cnt[22] ? _GEN_5528 : _GEN_5455; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_5666 = cnt[22] ? _GEN_5529 : _GEN_5456; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_5667 = cnt[22] ? _GEN_5530 : _GEN_5457; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_5668 = cnt[22] ? _GEN_5531 : _GEN_5458; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5669 = cnt[22] ? _GEN_5532 : _GEN_5459; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5670 = cnt[22] ? _GEN_5533 : _GEN_5460; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5671 = cnt[22] ? _GEN_5534 : _GEN_5461; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5672 = cnt[22] ? _GEN_5535 : _GEN_5462; // @[NulCtrlMP.scala 843:29]
  wire [128:0] _GEN_5673 = cnt[22] ? _GEN_5600 : _GEN_5463; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5674 = cnt[22] ? _GEN_5601 : _GEN_5464; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5675 = cnt[22] ? _GEN_5602 : _GEN_5465; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5676 = cnt[22] ? _GEN_5603 : _GEN_5466; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5677 = cnt[22] ? _GEN_5604 : _GEN_5467; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5678 = cnt[22] ? _GEN_5605 : _GEN_5468; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5679 = cnt[22] ? _GEN_5606 : _GEN_5469; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5680 = cnt[22] ? _GEN_5607 : _GEN_5470; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5681 = cnt[22] ? _GEN_5608 : _GEN_5471; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5682 = cnt[22] ? _GEN_5609 : _GEN_5472; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5683 = cnt[22] ? _GEN_5610 : _GEN_5473; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5684 = cnt[22] ? _GEN_5611 : _GEN_5474; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5685 = cnt[22] ? _GEN_5612 : _GEN_5475; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5686 = cnt[22] ? _GEN_5613 : _GEN_5476; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5687 = cnt[22] ? _GEN_5614 : _GEN_5477; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5688 = cnt[22] ? _GEN_5615 : _GEN_5478; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5689 = cnt[22] ? _GEN_5616 : _GEN_5479; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5690 = cnt[22] ? _GEN_5617 : _GEN_5480; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5691 = cnt[22] ? _GEN_5618 : _GEN_5481; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5692 = cnt[22] ? _GEN_5619 : _GEN_5482; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5693 = cnt[22] ? _GEN_5620 : _GEN_5483; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5694 = cnt[22] ? _GEN_5621 : _GEN_5484; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5695 = cnt[22] ? _GEN_5622 : _GEN_5485; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5696 = cnt[22] ? _GEN_5623 : _GEN_5486; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5697 = cnt[22] ? _GEN_5624 : _GEN_5487; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5698 = cnt[22] ? _GEN_5625 : _GEN_5488; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5699 = cnt[22] ? _GEN_5626 : _GEN_5489; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5700 = cnt[22] ? _GEN_5627 : _GEN_5490; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5701 = cnt[22] ? _GEN_5628 : _GEN_5491; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5702 = cnt[22] ? _GEN_5629 : _GEN_5492; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5703 = cnt[22] ? _GEN_5630 : _GEN_5493; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5704 = cnt[22] ? _GEN_5631 : _GEN_5494; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5705 = cnt[22] ? _GEN_5632 : _GEN_5495; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5706 = cnt[22] ? _GEN_5633 : _GEN_5496; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5707 = cnt[22] ? _GEN_5634 : _GEN_5497; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5708 = cnt[22] ? _GEN_5635 : _GEN_5498; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5709 = cnt[22] ? _GEN_5636 : _GEN_5499; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5710 = cnt[22] ? _GEN_5637 : _GEN_5500; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5711 = cnt[22] ? _GEN_5638 : _GEN_5501; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5712 = cnt[22] ? _GEN_5639 : _GEN_5502; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5713 = cnt[22] ? _GEN_5640 : _GEN_5503; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5714 = cnt[22] ? _GEN_5641 : _GEN_5504; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5715 = cnt[22] ? _GEN_5642 : _GEN_5505; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5716 = cnt[22] ? _GEN_5643 : _GEN_5506; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5717 = cnt[22] ? _GEN_5644 : _GEN_5507; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5718 = cnt[22] ? _GEN_5645 : _GEN_5508; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5719 = cnt[22] ? _GEN_5646 : _GEN_5509; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5720 = cnt[22] ? _GEN_5647 : _GEN_5510; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5721 = cnt[22] ? _GEN_5648 : _GEN_5511; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5722 = cnt[22] ? _GEN_5649 : _GEN_5512; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5723 = cnt[22] ? _GEN_5650 : _GEN_5513; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5724 = cnt[22] ? _GEN_5651 : _GEN_5514; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5725 = cnt[22] ? _GEN_5652 : _GEN_5515; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5726 = cnt[22] ? _GEN_5653 : _GEN_5516; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5727 = cnt[22] ? _GEN_5654 : _GEN_5517; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5728 = cnt[22] ? _GEN_5655 : _GEN_5518; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5729 = cnt[22] ? _GEN_5656 : _GEN_5519; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5730 = cnt[22] ? _GEN_5657 : _GEN_5520; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5731 = cnt[22] ? _GEN_5658 : _GEN_5521; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5732 = cnt[22] ? _GEN_5659 : _GEN_5522; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5733 = cnt[22] ? _GEN_5660 : _GEN_5523; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5734 = cnt[22] ? _GEN_5661 : _GEN_5524; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5735 = cnt[22] ? _GEN_5662 : _GEN_5525; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5736 = cnt[22] ? _GEN_5663 : _GEN_5526; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5737 = cnt[22] ? _GEN_5664 : _GEN_5527; // @[NulCtrlMP.scala 843:29]
  wire [8:0] _T_492 = pgbuf_cpu_pos[11:3] + 9'h2; // @[NulCtrlMP.scala 843:77]
  wire  _GEN_5738 = _GEN_145 | _GEN_5665; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5739 = _GEN_146 | _GEN_5666; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5740 = _GEN_147 | _GEN_5667; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5741 = _GEN_148 | _GEN_5668; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5742 = 2'h0 == opidx ? 5'h8 : _GEN_5669; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5743 = 2'h1 == opidx ? 5'h8 : _GEN_5670; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5744 = 2'h2 == opidx ? 5'h8 : _GEN_5671; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5745 = 2'h3 == opidx ? 5'h8 : _GEN_5672; // @[NulCtrlMP.scala 352:{28,28}]
  wire [63:0] _GEN_5746 = 6'h0 == _T_492[5:0] ? _GEN_1349 : _GEN_5674; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5747 = 6'h1 == _T_492[5:0] ? _GEN_1349 : _GEN_5675; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5748 = 6'h2 == _T_492[5:0] ? _GEN_1349 : _GEN_5676; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5749 = 6'h3 == _T_492[5:0] ? _GEN_1349 : _GEN_5677; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5750 = 6'h4 == _T_492[5:0] ? _GEN_1349 : _GEN_5678; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5751 = 6'h5 == _T_492[5:0] ? _GEN_1349 : _GEN_5679; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5752 = 6'h6 == _T_492[5:0] ? _GEN_1349 : _GEN_5680; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5753 = 6'h7 == _T_492[5:0] ? _GEN_1349 : _GEN_5681; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5754 = 6'h8 == _T_492[5:0] ? _GEN_1349 : _GEN_5682; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5755 = 6'h9 == _T_492[5:0] ? _GEN_1349 : _GEN_5683; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5756 = 6'ha == _T_492[5:0] ? _GEN_1349 : _GEN_5684; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5757 = 6'hb == _T_492[5:0] ? _GEN_1349 : _GEN_5685; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5758 = 6'hc == _T_492[5:0] ? _GEN_1349 : _GEN_5686; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5759 = 6'hd == _T_492[5:0] ? _GEN_1349 : _GEN_5687; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5760 = 6'he == _T_492[5:0] ? _GEN_1349 : _GEN_5688; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5761 = 6'hf == _T_492[5:0] ? _GEN_1349 : _GEN_5689; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5762 = 6'h10 == _T_492[5:0] ? _GEN_1349 : _GEN_5690; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5763 = 6'h11 == _T_492[5:0] ? _GEN_1349 : _GEN_5691; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5764 = 6'h12 == _T_492[5:0] ? _GEN_1349 : _GEN_5692; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5765 = 6'h13 == _T_492[5:0] ? _GEN_1349 : _GEN_5693; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5766 = 6'h14 == _T_492[5:0] ? _GEN_1349 : _GEN_5694; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5767 = 6'h15 == _T_492[5:0] ? _GEN_1349 : _GEN_5695; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5768 = 6'h16 == _T_492[5:0] ? _GEN_1349 : _GEN_5696; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5769 = 6'h17 == _T_492[5:0] ? _GEN_1349 : _GEN_5697; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5770 = 6'h18 == _T_492[5:0] ? _GEN_1349 : _GEN_5698; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5771 = 6'h19 == _T_492[5:0] ? _GEN_1349 : _GEN_5699; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5772 = 6'h1a == _T_492[5:0] ? _GEN_1349 : _GEN_5700; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5773 = 6'h1b == _T_492[5:0] ? _GEN_1349 : _GEN_5701; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5774 = 6'h1c == _T_492[5:0] ? _GEN_1349 : _GEN_5702; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5775 = 6'h1d == _T_492[5:0] ? _GEN_1349 : _GEN_5703; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5776 = 6'h1e == _T_492[5:0] ? _GEN_1349 : _GEN_5704; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5777 = 6'h1f == _T_492[5:0] ? _GEN_1349 : _GEN_5705; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5778 = 6'h20 == _T_492[5:0] ? _GEN_1349 : _GEN_5706; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5779 = 6'h21 == _T_492[5:0] ? _GEN_1349 : _GEN_5707; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5780 = 6'h22 == _T_492[5:0] ? _GEN_1349 : _GEN_5708; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5781 = 6'h23 == _T_492[5:0] ? _GEN_1349 : _GEN_5709; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5782 = 6'h24 == _T_492[5:0] ? _GEN_1349 : _GEN_5710; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5783 = 6'h25 == _T_492[5:0] ? _GEN_1349 : _GEN_5711; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5784 = 6'h26 == _T_492[5:0] ? _GEN_1349 : _GEN_5712; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5785 = 6'h27 == _T_492[5:0] ? _GEN_1349 : _GEN_5713; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5786 = 6'h28 == _T_492[5:0] ? _GEN_1349 : _GEN_5714; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5787 = 6'h29 == _T_492[5:0] ? _GEN_1349 : _GEN_5715; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5788 = 6'h2a == _T_492[5:0] ? _GEN_1349 : _GEN_5716; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5789 = 6'h2b == _T_492[5:0] ? _GEN_1349 : _GEN_5717; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5790 = 6'h2c == _T_492[5:0] ? _GEN_1349 : _GEN_5718; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5791 = 6'h2d == _T_492[5:0] ? _GEN_1349 : _GEN_5719; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5792 = 6'h2e == _T_492[5:0] ? _GEN_1349 : _GEN_5720; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5793 = 6'h2f == _T_492[5:0] ? _GEN_1349 : _GEN_5721; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5794 = 6'h30 == _T_492[5:0] ? _GEN_1349 : _GEN_5722; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5795 = 6'h31 == _T_492[5:0] ? _GEN_1349 : _GEN_5723; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5796 = 6'h32 == _T_492[5:0] ? _GEN_1349 : _GEN_5724; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5797 = 6'h33 == _T_492[5:0] ? _GEN_1349 : _GEN_5725; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5798 = 6'h34 == _T_492[5:0] ? _GEN_1349 : _GEN_5726; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5799 = 6'h35 == _T_492[5:0] ? _GEN_1349 : _GEN_5727; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5800 = 6'h36 == _T_492[5:0] ? _GEN_1349 : _GEN_5728; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5801 = 6'h37 == _T_492[5:0] ? _GEN_1349 : _GEN_5729; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5802 = 6'h38 == _T_492[5:0] ? _GEN_1349 : _GEN_5730; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5803 = 6'h39 == _T_492[5:0] ? _GEN_1349 : _GEN_5731; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5804 = 6'h3a == _T_492[5:0] ? _GEN_1349 : _GEN_5732; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5805 = 6'h3b == _T_492[5:0] ? _GEN_1349 : _GEN_5733; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5806 = 6'h3c == _T_492[5:0] ? _GEN_1349 : _GEN_5734; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5807 = 6'h3d == _T_492[5:0] ? _GEN_1349 : _GEN_5735; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5808 = 6'h3e == _T_492[5:0] ? _GEN_1349 : _GEN_5736; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5809 = 6'h3f == _T_492[5:0] ? _GEN_1349 : _GEN_5737; // @[NulCtrlMP.scala 355:{17,17}]
  wire [128:0] _GEN_5810 = _T_122 ? _cnt_T : _GEN_5673; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_5811 = _T_122 ? _GEN_5746 : _GEN_5674; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5812 = _T_122 ? _GEN_5747 : _GEN_5675; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5813 = _T_122 ? _GEN_5748 : _GEN_5676; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5814 = _T_122 ? _GEN_5749 : _GEN_5677; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5815 = _T_122 ? _GEN_5750 : _GEN_5678; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5816 = _T_122 ? _GEN_5751 : _GEN_5679; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5817 = _T_122 ? _GEN_5752 : _GEN_5680; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5818 = _T_122 ? _GEN_5753 : _GEN_5681; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5819 = _T_122 ? _GEN_5754 : _GEN_5682; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5820 = _T_122 ? _GEN_5755 : _GEN_5683; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5821 = _T_122 ? _GEN_5756 : _GEN_5684; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5822 = _T_122 ? _GEN_5757 : _GEN_5685; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5823 = _T_122 ? _GEN_5758 : _GEN_5686; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5824 = _T_122 ? _GEN_5759 : _GEN_5687; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5825 = _T_122 ? _GEN_5760 : _GEN_5688; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5826 = _T_122 ? _GEN_5761 : _GEN_5689; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5827 = _T_122 ? _GEN_5762 : _GEN_5690; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5828 = _T_122 ? _GEN_5763 : _GEN_5691; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5829 = _T_122 ? _GEN_5764 : _GEN_5692; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5830 = _T_122 ? _GEN_5765 : _GEN_5693; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5831 = _T_122 ? _GEN_5766 : _GEN_5694; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5832 = _T_122 ? _GEN_5767 : _GEN_5695; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5833 = _T_122 ? _GEN_5768 : _GEN_5696; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5834 = _T_122 ? _GEN_5769 : _GEN_5697; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5835 = _T_122 ? _GEN_5770 : _GEN_5698; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5836 = _T_122 ? _GEN_5771 : _GEN_5699; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5837 = _T_122 ? _GEN_5772 : _GEN_5700; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5838 = _T_122 ? _GEN_5773 : _GEN_5701; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5839 = _T_122 ? _GEN_5774 : _GEN_5702; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5840 = _T_122 ? _GEN_5775 : _GEN_5703; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5841 = _T_122 ? _GEN_5776 : _GEN_5704; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5842 = _T_122 ? _GEN_5777 : _GEN_5705; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5843 = _T_122 ? _GEN_5778 : _GEN_5706; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5844 = _T_122 ? _GEN_5779 : _GEN_5707; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5845 = _T_122 ? _GEN_5780 : _GEN_5708; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5846 = _T_122 ? _GEN_5781 : _GEN_5709; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5847 = _T_122 ? _GEN_5782 : _GEN_5710; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5848 = _T_122 ? _GEN_5783 : _GEN_5711; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5849 = _T_122 ? _GEN_5784 : _GEN_5712; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5850 = _T_122 ? _GEN_5785 : _GEN_5713; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5851 = _T_122 ? _GEN_5786 : _GEN_5714; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5852 = _T_122 ? _GEN_5787 : _GEN_5715; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5853 = _T_122 ? _GEN_5788 : _GEN_5716; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5854 = _T_122 ? _GEN_5789 : _GEN_5717; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5855 = _T_122 ? _GEN_5790 : _GEN_5718; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5856 = _T_122 ? _GEN_5791 : _GEN_5719; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5857 = _T_122 ? _GEN_5792 : _GEN_5720; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5858 = _T_122 ? _GEN_5793 : _GEN_5721; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5859 = _T_122 ? _GEN_5794 : _GEN_5722; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5860 = _T_122 ? _GEN_5795 : _GEN_5723; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5861 = _T_122 ? _GEN_5796 : _GEN_5724; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5862 = _T_122 ? _GEN_5797 : _GEN_5725; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5863 = _T_122 ? _GEN_5798 : _GEN_5726; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5864 = _T_122 ? _GEN_5799 : _GEN_5727; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5865 = _T_122 ? _GEN_5800 : _GEN_5728; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5866 = _T_122 ? _GEN_5801 : _GEN_5729; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5867 = _T_122 ? _GEN_5802 : _GEN_5730; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5868 = _T_122 ? _GEN_5803 : _GEN_5731; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5869 = _T_122 ? _GEN_5804 : _GEN_5732; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5870 = _T_122 ? _GEN_5805 : _GEN_5733; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5871 = _T_122 ? _GEN_5806 : _GEN_5734; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5872 = _T_122 ? _GEN_5807 : _GEN_5735; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5873 = _T_122 ? _GEN_5808 : _GEN_5736; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_5874 = _T_122 ? _GEN_5809 : _GEN_5737; // @[NulCtrlMP.scala 353:36]
  wire  _GEN_5875 = cnt[23] ? _GEN_5738 : _GEN_5665; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_5876 = cnt[23] ? _GEN_5739 : _GEN_5666; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_5877 = cnt[23] ? _GEN_5740 : _GEN_5667; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_5878 = cnt[23] ? _GEN_5741 : _GEN_5668; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5879 = cnt[23] ? _GEN_5742 : _GEN_5669; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5880 = cnt[23] ? _GEN_5743 : _GEN_5670; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5881 = cnt[23] ? _GEN_5744 : _GEN_5671; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_5882 = cnt[23] ? _GEN_5745 : _GEN_5672; // @[NulCtrlMP.scala 843:29]
  wire [128:0] _GEN_5883 = cnt[23] ? _GEN_5810 : _GEN_5673; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5884 = cnt[23] ? _GEN_5811 : _GEN_5674; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5885 = cnt[23] ? _GEN_5812 : _GEN_5675; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5886 = cnt[23] ? _GEN_5813 : _GEN_5676; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5887 = cnt[23] ? _GEN_5814 : _GEN_5677; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5888 = cnt[23] ? _GEN_5815 : _GEN_5678; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5889 = cnt[23] ? _GEN_5816 : _GEN_5679; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5890 = cnt[23] ? _GEN_5817 : _GEN_5680; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5891 = cnt[23] ? _GEN_5818 : _GEN_5681; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5892 = cnt[23] ? _GEN_5819 : _GEN_5682; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5893 = cnt[23] ? _GEN_5820 : _GEN_5683; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5894 = cnt[23] ? _GEN_5821 : _GEN_5684; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5895 = cnt[23] ? _GEN_5822 : _GEN_5685; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5896 = cnt[23] ? _GEN_5823 : _GEN_5686; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5897 = cnt[23] ? _GEN_5824 : _GEN_5687; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5898 = cnt[23] ? _GEN_5825 : _GEN_5688; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5899 = cnt[23] ? _GEN_5826 : _GEN_5689; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5900 = cnt[23] ? _GEN_5827 : _GEN_5690; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5901 = cnt[23] ? _GEN_5828 : _GEN_5691; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5902 = cnt[23] ? _GEN_5829 : _GEN_5692; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5903 = cnt[23] ? _GEN_5830 : _GEN_5693; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5904 = cnt[23] ? _GEN_5831 : _GEN_5694; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5905 = cnt[23] ? _GEN_5832 : _GEN_5695; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5906 = cnt[23] ? _GEN_5833 : _GEN_5696; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5907 = cnt[23] ? _GEN_5834 : _GEN_5697; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5908 = cnt[23] ? _GEN_5835 : _GEN_5698; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5909 = cnt[23] ? _GEN_5836 : _GEN_5699; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5910 = cnt[23] ? _GEN_5837 : _GEN_5700; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5911 = cnt[23] ? _GEN_5838 : _GEN_5701; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5912 = cnt[23] ? _GEN_5839 : _GEN_5702; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5913 = cnt[23] ? _GEN_5840 : _GEN_5703; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5914 = cnt[23] ? _GEN_5841 : _GEN_5704; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5915 = cnt[23] ? _GEN_5842 : _GEN_5705; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5916 = cnt[23] ? _GEN_5843 : _GEN_5706; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5917 = cnt[23] ? _GEN_5844 : _GEN_5707; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5918 = cnt[23] ? _GEN_5845 : _GEN_5708; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5919 = cnt[23] ? _GEN_5846 : _GEN_5709; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5920 = cnt[23] ? _GEN_5847 : _GEN_5710; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5921 = cnt[23] ? _GEN_5848 : _GEN_5711; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5922 = cnt[23] ? _GEN_5849 : _GEN_5712; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5923 = cnt[23] ? _GEN_5850 : _GEN_5713; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5924 = cnt[23] ? _GEN_5851 : _GEN_5714; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5925 = cnt[23] ? _GEN_5852 : _GEN_5715; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5926 = cnt[23] ? _GEN_5853 : _GEN_5716; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5927 = cnt[23] ? _GEN_5854 : _GEN_5717; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5928 = cnt[23] ? _GEN_5855 : _GEN_5718; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5929 = cnt[23] ? _GEN_5856 : _GEN_5719; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5930 = cnt[23] ? _GEN_5857 : _GEN_5720; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5931 = cnt[23] ? _GEN_5858 : _GEN_5721; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5932 = cnt[23] ? _GEN_5859 : _GEN_5722; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5933 = cnt[23] ? _GEN_5860 : _GEN_5723; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5934 = cnt[23] ? _GEN_5861 : _GEN_5724; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5935 = cnt[23] ? _GEN_5862 : _GEN_5725; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5936 = cnt[23] ? _GEN_5863 : _GEN_5726; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5937 = cnt[23] ? _GEN_5864 : _GEN_5727; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5938 = cnt[23] ? _GEN_5865 : _GEN_5728; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5939 = cnt[23] ? _GEN_5866 : _GEN_5729; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5940 = cnt[23] ? _GEN_5867 : _GEN_5730; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5941 = cnt[23] ? _GEN_5868 : _GEN_5731; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5942 = cnt[23] ? _GEN_5869 : _GEN_5732; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5943 = cnt[23] ? _GEN_5870 : _GEN_5733; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5944 = cnt[23] ? _GEN_5871 : _GEN_5734; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5945 = cnt[23] ? _GEN_5872 : _GEN_5735; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5946 = cnt[23] ? _GEN_5873 : _GEN_5736; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_5947 = cnt[23] ? _GEN_5874 : _GEN_5737; // @[NulCtrlMP.scala 843:29]
  wire [8:0] _T_498 = pgbuf_cpu_pos[11:3] + 9'h3; // @[NulCtrlMP.scala 843:77]
  wire  _GEN_5948 = _GEN_145 | _GEN_5875; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5949 = _GEN_146 | _GEN_5876; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5950 = _GEN_147 | _GEN_5877; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_5951 = _GEN_148 | _GEN_5878; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_5952 = 2'h0 == opidx ? 5'h9 : _GEN_5879; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5953 = 2'h1 == opidx ? 5'h9 : _GEN_5880; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5954 = 2'h2 == opidx ? 5'h9 : _GEN_5881; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_5955 = 2'h3 == opidx ? 5'h9 : _GEN_5882; // @[NulCtrlMP.scala 352:{28,28}]
  wire [63:0] _GEN_5956 = 6'h0 == _T_498[5:0] ? _GEN_1349 : _GEN_5884; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5957 = 6'h1 == _T_498[5:0] ? _GEN_1349 : _GEN_5885; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5958 = 6'h2 == _T_498[5:0] ? _GEN_1349 : _GEN_5886; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5959 = 6'h3 == _T_498[5:0] ? _GEN_1349 : _GEN_5887; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5960 = 6'h4 == _T_498[5:0] ? _GEN_1349 : _GEN_5888; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5961 = 6'h5 == _T_498[5:0] ? _GEN_1349 : _GEN_5889; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5962 = 6'h6 == _T_498[5:0] ? _GEN_1349 : _GEN_5890; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5963 = 6'h7 == _T_498[5:0] ? _GEN_1349 : _GEN_5891; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5964 = 6'h8 == _T_498[5:0] ? _GEN_1349 : _GEN_5892; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5965 = 6'h9 == _T_498[5:0] ? _GEN_1349 : _GEN_5893; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5966 = 6'ha == _T_498[5:0] ? _GEN_1349 : _GEN_5894; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5967 = 6'hb == _T_498[5:0] ? _GEN_1349 : _GEN_5895; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5968 = 6'hc == _T_498[5:0] ? _GEN_1349 : _GEN_5896; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5969 = 6'hd == _T_498[5:0] ? _GEN_1349 : _GEN_5897; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5970 = 6'he == _T_498[5:0] ? _GEN_1349 : _GEN_5898; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5971 = 6'hf == _T_498[5:0] ? _GEN_1349 : _GEN_5899; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5972 = 6'h10 == _T_498[5:0] ? _GEN_1349 : _GEN_5900; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5973 = 6'h11 == _T_498[5:0] ? _GEN_1349 : _GEN_5901; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5974 = 6'h12 == _T_498[5:0] ? _GEN_1349 : _GEN_5902; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5975 = 6'h13 == _T_498[5:0] ? _GEN_1349 : _GEN_5903; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5976 = 6'h14 == _T_498[5:0] ? _GEN_1349 : _GEN_5904; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5977 = 6'h15 == _T_498[5:0] ? _GEN_1349 : _GEN_5905; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5978 = 6'h16 == _T_498[5:0] ? _GEN_1349 : _GEN_5906; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5979 = 6'h17 == _T_498[5:0] ? _GEN_1349 : _GEN_5907; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5980 = 6'h18 == _T_498[5:0] ? _GEN_1349 : _GEN_5908; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5981 = 6'h19 == _T_498[5:0] ? _GEN_1349 : _GEN_5909; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5982 = 6'h1a == _T_498[5:0] ? _GEN_1349 : _GEN_5910; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5983 = 6'h1b == _T_498[5:0] ? _GEN_1349 : _GEN_5911; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5984 = 6'h1c == _T_498[5:0] ? _GEN_1349 : _GEN_5912; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5985 = 6'h1d == _T_498[5:0] ? _GEN_1349 : _GEN_5913; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5986 = 6'h1e == _T_498[5:0] ? _GEN_1349 : _GEN_5914; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5987 = 6'h1f == _T_498[5:0] ? _GEN_1349 : _GEN_5915; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5988 = 6'h20 == _T_498[5:0] ? _GEN_1349 : _GEN_5916; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5989 = 6'h21 == _T_498[5:0] ? _GEN_1349 : _GEN_5917; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5990 = 6'h22 == _T_498[5:0] ? _GEN_1349 : _GEN_5918; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5991 = 6'h23 == _T_498[5:0] ? _GEN_1349 : _GEN_5919; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5992 = 6'h24 == _T_498[5:0] ? _GEN_1349 : _GEN_5920; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5993 = 6'h25 == _T_498[5:0] ? _GEN_1349 : _GEN_5921; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5994 = 6'h26 == _T_498[5:0] ? _GEN_1349 : _GEN_5922; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5995 = 6'h27 == _T_498[5:0] ? _GEN_1349 : _GEN_5923; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5996 = 6'h28 == _T_498[5:0] ? _GEN_1349 : _GEN_5924; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5997 = 6'h29 == _T_498[5:0] ? _GEN_1349 : _GEN_5925; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5998 = 6'h2a == _T_498[5:0] ? _GEN_1349 : _GEN_5926; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_5999 = 6'h2b == _T_498[5:0] ? _GEN_1349 : _GEN_5927; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6000 = 6'h2c == _T_498[5:0] ? _GEN_1349 : _GEN_5928; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6001 = 6'h2d == _T_498[5:0] ? _GEN_1349 : _GEN_5929; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6002 = 6'h2e == _T_498[5:0] ? _GEN_1349 : _GEN_5930; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6003 = 6'h2f == _T_498[5:0] ? _GEN_1349 : _GEN_5931; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6004 = 6'h30 == _T_498[5:0] ? _GEN_1349 : _GEN_5932; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6005 = 6'h31 == _T_498[5:0] ? _GEN_1349 : _GEN_5933; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6006 = 6'h32 == _T_498[5:0] ? _GEN_1349 : _GEN_5934; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6007 = 6'h33 == _T_498[5:0] ? _GEN_1349 : _GEN_5935; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6008 = 6'h34 == _T_498[5:0] ? _GEN_1349 : _GEN_5936; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6009 = 6'h35 == _T_498[5:0] ? _GEN_1349 : _GEN_5937; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6010 = 6'h36 == _T_498[5:0] ? _GEN_1349 : _GEN_5938; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6011 = 6'h37 == _T_498[5:0] ? _GEN_1349 : _GEN_5939; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6012 = 6'h38 == _T_498[5:0] ? _GEN_1349 : _GEN_5940; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6013 = 6'h39 == _T_498[5:0] ? _GEN_1349 : _GEN_5941; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6014 = 6'h3a == _T_498[5:0] ? _GEN_1349 : _GEN_5942; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6015 = 6'h3b == _T_498[5:0] ? _GEN_1349 : _GEN_5943; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6016 = 6'h3c == _T_498[5:0] ? _GEN_1349 : _GEN_5944; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6017 = 6'h3d == _T_498[5:0] ? _GEN_1349 : _GEN_5945; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6018 = 6'h3e == _T_498[5:0] ? _GEN_1349 : _GEN_5946; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6019 = 6'h3f == _T_498[5:0] ? _GEN_1349 : _GEN_5947; // @[NulCtrlMP.scala 355:{17,17}]
  wire [128:0] _GEN_6020 = _T_122 ? _cnt_T : _GEN_5883; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_6021 = _T_122 ? _GEN_5956 : _GEN_5884; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6022 = _T_122 ? _GEN_5957 : _GEN_5885; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6023 = _T_122 ? _GEN_5958 : _GEN_5886; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6024 = _T_122 ? _GEN_5959 : _GEN_5887; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6025 = _T_122 ? _GEN_5960 : _GEN_5888; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6026 = _T_122 ? _GEN_5961 : _GEN_5889; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6027 = _T_122 ? _GEN_5962 : _GEN_5890; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6028 = _T_122 ? _GEN_5963 : _GEN_5891; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6029 = _T_122 ? _GEN_5964 : _GEN_5892; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6030 = _T_122 ? _GEN_5965 : _GEN_5893; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6031 = _T_122 ? _GEN_5966 : _GEN_5894; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6032 = _T_122 ? _GEN_5967 : _GEN_5895; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6033 = _T_122 ? _GEN_5968 : _GEN_5896; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6034 = _T_122 ? _GEN_5969 : _GEN_5897; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6035 = _T_122 ? _GEN_5970 : _GEN_5898; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6036 = _T_122 ? _GEN_5971 : _GEN_5899; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6037 = _T_122 ? _GEN_5972 : _GEN_5900; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6038 = _T_122 ? _GEN_5973 : _GEN_5901; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6039 = _T_122 ? _GEN_5974 : _GEN_5902; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6040 = _T_122 ? _GEN_5975 : _GEN_5903; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6041 = _T_122 ? _GEN_5976 : _GEN_5904; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6042 = _T_122 ? _GEN_5977 : _GEN_5905; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6043 = _T_122 ? _GEN_5978 : _GEN_5906; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6044 = _T_122 ? _GEN_5979 : _GEN_5907; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6045 = _T_122 ? _GEN_5980 : _GEN_5908; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6046 = _T_122 ? _GEN_5981 : _GEN_5909; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6047 = _T_122 ? _GEN_5982 : _GEN_5910; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6048 = _T_122 ? _GEN_5983 : _GEN_5911; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6049 = _T_122 ? _GEN_5984 : _GEN_5912; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6050 = _T_122 ? _GEN_5985 : _GEN_5913; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6051 = _T_122 ? _GEN_5986 : _GEN_5914; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6052 = _T_122 ? _GEN_5987 : _GEN_5915; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6053 = _T_122 ? _GEN_5988 : _GEN_5916; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6054 = _T_122 ? _GEN_5989 : _GEN_5917; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6055 = _T_122 ? _GEN_5990 : _GEN_5918; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6056 = _T_122 ? _GEN_5991 : _GEN_5919; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6057 = _T_122 ? _GEN_5992 : _GEN_5920; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6058 = _T_122 ? _GEN_5993 : _GEN_5921; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6059 = _T_122 ? _GEN_5994 : _GEN_5922; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6060 = _T_122 ? _GEN_5995 : _GEN_5923; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6061 = _T_122 ? _GEN_5996 : _GEN_5924; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6062 = _T_122 ? _GEN_5997 : _GEN_5925; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6063 = _T_122 ? _GEN_5998 : _GEN_5926; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6064 = _T_122 ? _GEN_5999 : _GEN_5927; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6065 = _T_122 ? _GEN_6000 : _GEN_5928; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6066 = _T_122 ? _GEN_6001 : _GEN_5929; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6067 = _T_122 ? _GEN_6002 : _GEN_5930; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6068 = _T_122 ? _GEN_6003 : _GEN_5931; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6069 = _T_122 ? _GEN_6004 : _GEN_5932; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6070 = _T_122 ? _GEN_6005 : _GEN_5933; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6071 = _T_122 ? _GEN_6006 : _GEN_5934; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6072 = _T_122 ? _GEN_6007 : _GEN_5935; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6073 = _T_122 ? _GEN_6008 : _GEN_5936; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6074 = _T_122 ? _GEN_6009 : _GEN_5937; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6075 = _T_122 ? _GEN_6010 : _GEN_5938; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6076 = _T_122 ? _GEN_6011 : _GEN_5939; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6077 = _T_122 ? _GEN_6012 : _GEN_5940; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6078 = _T_122 ? _GEN_6013 : _GEN_5941; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6079 = _T_122 ? _GEN_6014 : _GEN_5942; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6080 = _T_122 ? _GEN_6015 : _GEN_5943; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6081 = _T_122 ? _GEN_6016 : _GEN_5944; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6082 = _T_122 ? _GEN_6017 : _GEN_5945; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6083 = _T_122 ? _GEN_6018 : _GEN_5946; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6084 = _T_122 ? _GEN_6019 : _GEN_5947; // @[NulCtrlMP.scala 353:36]
  wire  _GEN_6085 = cnt[24] ? _GEN_5948 : _GEN_5875; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6086 = cnt[24] ? _GEN_5949 : _GEN_5876; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6087 = cnt[24] ? _GEN_5950 : _GEN_5877; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6088 = cnt[24] ? _GEN_5951 : _GEN_5878; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6089 = cnt[24] ? _GEN_5952 : _GEN_5879; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6090 = cnt[24] ? _GEN_5953 : _GEN_5880; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6091 = cnt[24] ? _GEN_5954 : _GEN_5881; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6092 = cnt[24] ? _GEN_5955 : _GEN_5882; // @[NulCtrlMP.scala 843:29]
  wire [128:0] _GEN_6093 = cnt[24] ? _GEN_6020 : _GEN_5883; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6094 = cnt[24] ? _GEN_6021 : _GEN_5884; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6095 = cnt[24] ? _GEN_6022 : _GEN_5885; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6096 = cnt[24] ? _GEN_6023 : _GEN_5886; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6097 = cnt[24] ? _GEN_6024 : _GEN_5887; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6098 = cnt[24] ? _GEN_6025 : _GEN_5888; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6099 = cnt[24] ? _GEN_6026 : _GEN_5889; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6100 = cnt[24] ? _GEN_6027 : _GEN_5890; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6101 = cnt[24] ? _GEN_6028 : _GEN_5891; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6102 = cnt[24] ? _GEN_6029 : _GEN_5892; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6103 = cnt[24] ? _GEN_6030 : _GEN_5893; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6104 = cnt[24] ? _GEN_6031 : _GEN_5894; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6105 = cnt[24] ? _GEN_6032 : _GEN_5895; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6106 = cnt[24] ? _GEN_6033 : _GEN_5896; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6107 = cnt[24] ? _GEN_6034 : _GEN_5897; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6108 = cnt[24] ? _GEN_6035 : _GEN_5898; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6109 = cnt[24] ? _GEN_6036 : _GEN_5899; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6110 = cnt[24] ? _GEN_6037 : _GEN_5900; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6111 = cnt[24] ? _GEN_6038 : _GEN_5901; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6112 = cnt[24] ? _GEN_6039 : _GEN_5902; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6113 = cnt[24] ? _GEN_6040 : _GEN_5903; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6114 = cnt[24] ? _GEN_6041 : _GEN_5904; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6115 = cnt[24] ? _GEN_6042 : _GEN_5905; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6116 = cnt[24] ? _GEN_6043 : _GEN_5906; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6117 = cnt[24] ? _GEN_6044 : _GEN_5907; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6118 = cnt[24] ? _GEN_6045 : _GEN_5908; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6119 = cnt[24] ? _GEN_6046 : _GEN_5909; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6120 = cnt[24] ? _GEN_6047 : _GEN_5910; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6121 = cnt[24] ? _GEN_6048 : _GEN_5911; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6122 = cnt[24] ? _GEN_6049 : _GEN_5912; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6123 = cnt[24] ? _GEN_6050 : _GEN_5913; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6124 = cnt[24] ? _GEN_6051 : _GEN_5914; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6125 = cnt[24] ? _GEN_6052 : _GEN_5915; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6126 = cnt[24] ? _GEN_6053 : _GEN_5916; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6127 = cnt[24] ? _GEN_6054 : _GEN_5917; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6128 = cnt[24] ? _GEN_6055 : _GEN_5918; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6129 = cnt[24] ? _GEN_6056 : _GEN_5919; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6130 = cnt[24] ? _GEN_6057 : _GEN_5920; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6131 = cnt[24] ? _GEN_6058 : _GEN_5921; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6132 = cnt[24] ? _GEN_6059 : _GEN_5922; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6133 = cnt[24] ? _GEN_6060 : _GEN_5923; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6134 = cnt[24] ? _GEN_6061 : _GEN_5924; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6135 = cnt[24] ? _GEN_6062 : _GEN_5925; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6136 = cnt[24] ? _GEN_6063 : _GEN_5926; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6137 = cnt[24] ? _GEN_6064 : _GEN_5927; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6138 = cnt[24] ? _GEN_6065 : _GEN_5928; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6139 = cnt[24] ? _GEN_6066 : _GEN_5929; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6140 = cnt[24] ? _GEN_6067 : _GEN_5930; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6141 = cnt[24] ? _GEN_6068 : _GEN_5931; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6142 = cnt[24] ? _GEN_6069 : _GEN_5932; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6143 = cnt[24] ? _GEN_6070 : _GEN_5933; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6144 = cnt[24] ? _GEN_6071 : _GEN_5934; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6145 = cnt[24] ? _GEN_6072 : _GEN_5935; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6146 = cnt[24] ? _GEN_6073 : _GEN_5936; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6147 = cnt[24] ? _GEN_6074 : _GEN_5937; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6148 = cnt[24] ? _GEN_6075 : _GEN_5938; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6149 = cnt[24] ? _GEN_6076 : _GEN_5939; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6150 = cnt[24] ? _GEN_6077 : _GEN_5940; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6151 = cnt[24] ? _GEN_6078 : _GEN_5941; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6152 = cnt[24] ? _GEN_6079 : _GEN_5942; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6153 = cnt[24] ? _GEN_6080 : _GEN_5943; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6154 = cnt[24] ? _GEN_6081 : _GEN_5944; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6155 = cnt[24] ? _GEN_6082 : _GEN_5945; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6156 = cnt[24] ? _GEN_6083 : _GEN_5946; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6157 = cnt[24] ? _GEN_6084 : _GEN_5947; // @[NulCtrlMP.scala 843:29]
  wire [8:0] _T_504 = pgbuf_cpu_pos[11:3] + 9'h4; // @[NulCtrlMP.scala 843:77]
  wire  _GEN_6158 = _GEN_145 | _GEN_6085; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6159 = _GEN_146 | _GEN_6086; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6160 = _GEN_147 | _GEN_6087; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6161 = _GEN_148 | _GEN_6088; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_6162 = 2'h0 == opidx ? 5'ha : _GEN_6089; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6163 = 2'h1 == opidx ? 5'ha : _GEN_6090; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6164 = 2'h2 == opidx ? 5'ha : _GEN_6091; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6165 = 2'h3 == opidx ? 5'ha : _GEN_6092; // @[NulCtrlMP.scala 352:{28,28}]
  wire [63:0] _GEN_6166 = 6'h0 == _T_504[5:0] ? _GEN_1349 : _GEN_6094; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6167 = 6'h1 == _T_504[5:0] ? _GEN_1349 : _GEN_6095; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6168 = 6'h2 == _T_504[5:0] ? _GEN_1349 : _GEN_6096; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6169 = 6'h3 == _T_504[5:0] ? _GEN_1349 : _GEN_6097; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6170 = 6'h4 == _T_504[5:0] ? _GEN_1349 : _GEN_6098; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6171 = 6'h5 == _T_504[5:0] ? _GEN_1349 : _GEN_6099; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6172 = 6'h6 == _T_504[5:0] ? _GEN_1349 : _GEN_6100; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6173 = 6'h7 == _T_504[5:0] ? _GEN_1349 : _GEN_6101; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6174 = 6'h8 == _T_504[5:0] ? _GEN_1349 : _GEN_6102; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6175 = 6'h9 == _T_504[5:0] ? _GEN_1349 : _GEN_6103; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6176 = 6'ha == _T_504[5:0] ? _GEN_1349 : _GEN_6104; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6177 = 6'hb == _T_504[5:0] ? _GEN_1349 : _GEN_6105; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6178 = 6'hc == _T_504[5:0] ? _GEN_1349 : _GEN_6106; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6179 = 6'hd == _T_504[5:0] ? _GEN_1349 : _GEN_6107; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6180 = 6'he == _T_504[5:0] ? _GEN_1349 : _GEN_6108; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6181 = 6'hf == _T_504[5:0] ? _GEN_1349 : _GEN_6109; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6182 = 6'h10 == _T_504[5:0] ? _GEN_1349 : _GEN_6110; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6183 = 6'h11 == _T_504[5:0] ? _GEN_1349 : _GEN_6111; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6184 = 6'h12 == _T_504[5:0] ? _GEN_1349 : _GEN_6112; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6185 = 6'h13 == _T_504[5:0] ? _GEN_1349 : _GEN_6113; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6186 = 6'h14 == _T_504[5:0] ? _GEN_1349 : _GEN_6114; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6187 = 6'h15 == _T_504[5:0] ? _GEN_1349 : _GEN_6115; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6188 = 6'h16 == _T_504[5:0] ? _GEN_1349 : _GEN_6116; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6189 = 6'h17 == _T_504[5:0] ? _GEN_1349 : _GEN_6117; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6190 = 6'h18 == _T_504[5:0] ? _GEN_1349 : _GEN_6118; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6191 = 6'h19 == _T_504[5:0] ? _GEN_1349 : _GEN_6119; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6192 = 6'h1a == _T_504[5:0] ? _GEN_1349 : _GEN_6120; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6193 = 6'h1b == _T_504[5:0] ? _GEN_1349 : _GEN_6121; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6194 = 6'h1c == _T_504[5:0] ? _GEN_1349 : _GEN_6122; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6195 = 6'h1d == _T_504[5:0] ? _GEN_1349 : _GEN_6123; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6196 = 6'h1e == _T_504[5:0] ? _GEN_1349 : _GEN_6124; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6197 = 6'h1f == _T_504[5:0] ? _GEN_1349 : _GEN_6125; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6198 = 6'h20 == _T_504[5:0] ? _GEN_1349 : _GEN_6126; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6199 = 6'h21 == _T_504[5:0] ? _GEN_1349 : _GEN_6127; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6200 = 6'h22 == _T_504[5:0] ? _GEN_1349 : _GEN_6128; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6201 = 6'h23 == _T_504[5:0] ? _GEN_1349 : _GEN_6129; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6202 = 6'h24 == _T_504[5:0] ? _GEN_1349 : _GEN_6130; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6203 = 6'h25 == _T_504[5:0] ? _GEN_1349 : _GEN_6131; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6204 = 6'h26 == _T_504[5:0] ? _GEN_1349 : _GEN_6132; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6205 = 6'h27 == _T_504[5:0] ? _GEN_1349 : _GEN_6133; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6206 = 6'h28 == _T_504[5:0] ? _GEN_1349 : _GEN_6134; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6207 = 6'h29 == _T_504[5:0] ? _GEN_1349 : _GEN_6135; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6208 = 6'h2a == _T_504[5:0] ? _GEN_1349 : _GEN_6136; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6209 = 6'h2b == _T_504[5:0] ? _GEN_1349 : _GEN_6137; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6210 = 6'h2c == _T_504[5:0] ? _GEN_1349 : _GEN_6138; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6211 = 6'h2d == _T_504[5:0] ? _GEN_1349 : _GEN_6139; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6212 = 6'h2e == _T_504[5:0] ? _GEN_1349 : _GEN_6140; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6213 = 6'h2f == _T_504[5:0] ? _GEN_1349 : _GEN_6141; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6214 = 6'h30 == _T_504[5:0] ? _GEN_1349 : _GEN_6142; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6215 = 6'h31 == _T_504[5:0] ? _GEN_1349 : _GEN_6143; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6216 = 6'h32 == _T_504[5:0] ? _GEN_1349 : _GEN_6144; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6217 = 6'h33 == _T_504[5:0] ? _GEN_1349 : _GEN_6145; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6218 = 6'h34 == _T_504[5:0] ? _GEN_1349 : _GEN_6146; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6219 = 6'h35 == _T_504[5:0] ? _GEN_1349 : _GEN_6147; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6220 = 6'h36 == _T_504[5:0] ? _GEN_1349 : _GEN_6148; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6221 = 6'h37 == _T_504[5:0] ? _GEN_1349 : _GEN_6149; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6222 = 6'h38 == _T_504[5:0] ? _GEN_1349 : _GEN_6150; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6223 = 6'h39 == _T_504[5:0] ? _GEN_1349 : _GEN_6151; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6224 = 6'h3a == _T_504[5:0] ? _GEN_1349 : _GEN_6152; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6225 = 6'h3b == _T_504[5:0] ? _GEN_1349 : _GEN_6153; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6226 = 6'h3c == _T_504[5:0] ? _GEN_1349 : _GEN_6154; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6227 = 6'h3d == _T_504[5:0] ? _GEN_1349 : _GEN_6155; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6228 = 6'h3e == _T_504[5:0] ? _GEN_1349 : _GEN_6156; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6229 = 6'h3f == _T_504[5:0] ? _GEN_1349 : _GEN_6157; // @[NulCtrlMP.scala 355:{17,17}]
  wire [128:0] _GEN_6230 = _T_122 ? _cnt_T : _GEN_6093; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_6231 = _T_122 ? _GEN_6166 : _GEN_6094; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6232 = _T_122 ? _GEN_6167 : _GEN_6095; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6233 = _T_122 ? _GEN_6168 : _GEN_6096; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6234 = _T_122 ? _GEN_6169 : _GEN_6097; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6235 = _T_122 ? _GEN_6170 : _GEN_6098; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6236 = _T_122 ? _GEN_6171 : _GEN_6099; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6237 = _T_122 ? _GEN_6172 : _GEN_6100; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6238 = _T_122 ? _GEN_6173 : _GEN_6101; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6239 = _T_122 ? _GEN_6174 : _GEN_6102; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6240 = _T_122 ? _GEN_6175 : _GEN_6103; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6241 = _T_122 ? _GEN_6176 : _GEN_6104; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6242 = _T_122 ? _GEN_6177 : _GEN_6105; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6243 = _T_122 ? _GEN_6178 : _GEN_6106; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6244 = _T_122 ? _GEN_6179 : _GEN_6107; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6245 = _T_122 ? _GEN_6180 : _GEN_6108; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6246 = _T_122 ? _GEN_6181 : _GEN_6109; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6247 = _T_122 ? _GEN_6182 : _GEN_6110; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6248 = _T_122 ? _GEN_6183 : _GEN_6111; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6249 = _T_122 ? _GEN_6184 : _GEN_6112; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6250 = _T_122 ? _GEN_6185 : _GEN_6113; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6251 = _T_122 ? _GEN_6186 : _GEN_6114; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6252 = _T_122 ? _GEN_6187 : _GEN_6115; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6253 = _T_122 ? _GEN_6188 : _GEN_6116; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6254 = _T_122 ? _GEN_6189 : _GEN_6117; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6255 = _T_122 ? _GEN_6190 : _GEN_6118; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6256 = _T_122 ? _GEN_6191 : _GEN_6119; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6257 = _T_122 ? _GEN_6192 : _GEN_6120; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6258 = _T_122 ? _GEN_6193 : _GEN_6121; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6259 = _T_122 ? _GEN_6194 : _GEN_6122; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6260 = _T_122 ? _GEN_6195 : _GEN_6123; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6261 = _T_122 ? _GEN_6196 : _GEN_6124; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6262 = _T_122 ? _GEN_6197 : _GEN_6125; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6263 = _T_122 ? _GEN_6198 : _GEN_6126; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6264 = _T_122 ? _GEN_6199 : _GEN_6127; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6265 = _T_122 ? _GEN_6200 : _GEN_6128; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6266 = _T_122 ? _GEN_6201 : _GEN_6129; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6267 = _T_122 ? _GEN_6202 : _GEN_6130; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6268 = _T_122 ? _GEN_6203 : _GEN_6131; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6269 = _T_122 ? _GEN_6204 : _GEN_6132; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6270 = _T_122 ? _GEN_6205 : _GEN_6133; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6271 = _T_122 ? _GEN_6206 : _GEN_6134; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6272 = _T_122 ? _GEN_6207 : _GEN_6135; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6273 = _T_122 ? _GEN_6208 : _GEN_6136; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6274 = _T_122 ? _GEN_6209 : _GEN_6137; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6275 = _T_122 ? _GEN_6210 : _GEN_6138; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6276 = _T_122 ? _GEN_6211 : _GEN_6139; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6277 = _T_122 ? _GEN_6212 : _GEN_6140; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6278 = _T_122 ? _GEN_6213 : _GEN_6141; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6279 = _T_122 ? _GEN_6214 : _GEN_6142; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6280 = _T_122 ? _GEN_6215 : _GEN_6143; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6281 = _T_122 ? _GEN_6216 : _GEN_6144; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6282 = _T_122 ? _GEN_6217 : _GEN_6145; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6283 = _T_122 ? _GEN_6218 : _GEN_6146; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6284 = _T_122 ? _GEN_6219 : _GEN_6147; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6285 = _T_122 ? _GEN_6220 : _GEN_6148; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6286 = _T_122 ? _GEN_6221 : _GEN_6149; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6287 = _T_122 ? _GEN_6222 : _GEN_6150; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6288 = _T_122 ? _GEN_6223 : _GEN_6151; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6289 = _T_122 ? _GEN_6224 : _GEN_6152; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6290 = _T_122 ? _GEN_6225 : _GEN_6153; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6291 = _T_122 ? _GEN_6226 : _GEN_6154; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6292 = _T_122 ? _GEN_6227 : _GEN_6155; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6293 = _T_122 ? _GEN_6228 : _GEN_6156; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6294 = _T_122 ? _GEN_6229 : _GEN_6157; // @[NulCtrlMP.scala 353:36]
  wire  _GEN_6295 = cnt[25] ? _GEN_6158 : _GEN_6085; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6296 = cnt[25] ? _GEN_6159 : _GEN_6086; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6297 = cnt[25] ? _GEN_6160 : _GEN_6087; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6298 = cnt[25] ? _GEN_6161 : _GEN_6088; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6299 = cnt[25] ? _GEN_6162 : _GEN_6089; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6300 = cnt[25] ? _GEN_6163 : _GEN_6090; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6301 = cnt[25] ? _GEN_6164 : _GEN_6091; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6302 = cnt[25] ? _GEN_6165 : _GEN_6092; // @[NulCtrlMP.scala 843:29]
  wire [128:0] _GEN_6303 = cnt[25] ? _GEN_6230 : _GEN_6093; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6304 = cnt[25] ? _GEN_6231 : _GEN_6094; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6305 = cnt[25] ? _GEN_6232 : _GEN_6095; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6306 = cnt[25] ? _GEN_6233 : _GEN_6096; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6307 = cnt[25] ? _GEN_6234 : _GEN_6097; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6308 = cnt[25] ? _GEN_6235 : _GEN_6098; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6309 = cnt[25] ? _GEN_6236 : _GEN_6099; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6310 = cnt[25] ? _GEN_6237 : _GEN_6100; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6311 = cnt[25] ? _GEN_6238 : _GEN_6101; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6312 = cnt[25] ? _GEN_6239 : _GEN_6102; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6313 = cnt[25] ? _GEN_6240 : _GEN_6103; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6314 = cnt[25] ? _GEN_6241 : _GEN_6104; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6315 = cnt[25] ? _GEN_6242 : _GEN_6105; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6316 = cnt[25] ? _GEN_6243 : _GEN_6106; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6317 = cnt[25] ? _GEN_6244 : _GEN_6107; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6318 = cnt[25] ? _GEN_6245 : _GEN_6108; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6319 = cnt[25] ? _GEN_6246 : _GEN_6109; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6320 = cnt[25] ? _GEN_6247 : _GEN_6110; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6321 = cnt[25] ? _GEN_6248 : _GEN_6111; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6322 = cnt[25] ? _GEN_6249 : _GEN_6112; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6323 = cnt[25] ? _GEN_6250 : _GEN_6113; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6324 = cnt[25] ? _GEN_6251 : _GEN_6114; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6325 = cnt[25] ? _GEN_6252 : _GEN_6115; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6326 = cnt[25] ? _GEN_6253 : _GEN_6116; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6327 = cnt[25] ? _GEN_6254 : _GEN_6117; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6328 = cnt[25] ? _GEN_6255 : _GEN_6118; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6329 = cnt[25] ? _GEN_6256 : _GEN_6119; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6330 = cnt[25] ? _GEN_6257 : _GEN_6120; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6331 = cnt[25] ? _GEN_6258 : _GEN_6121; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6332 = cnt[25] ? _GEN_6259 : _GEN_6122; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6333 = cnt[25] ? _GEN_6260 : _GEN_6123; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6334 = cnt[25] ? _GEN_6261 : _GEN_6124; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6335 = cnt[25] ? _GEN_6262 : _GEN_6125; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6336 = cnt[25] ? _GEN_6263 : _GEN_6126; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6337 = cnt[25] ? _GEN_6264 : _GEN_6127; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6338 = cnt[25] ? _GEN_6265 : _GEN_6128; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6339 = cnt[25] ? _GEN_6266 : _GEN_6129; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6340 = cnt[25] ? _GEN_6267 : _GEN_6130; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6341 = cnt[25] ? _GEN_6268 : _GEN_6131; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6342 = cnt[25] ? _GEN_6269 : _GEN_6132; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6343 = cnt[25] ? _GEN_6270 : _GEN_6133; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6344 = cnt[25] ? _GEN_6271 : _GEN_6134; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6345 = cnt[25] ? _GEN_6272 : _GEN_6135; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6346 = cnt[25] ? _GEN_6273 : _GEN_6136; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6347 = cnt[25] ? _GEN_6274 : _GEN_6137; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6348 = cnt[25] ? _GEN_6275 : _GEN_6138; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6349 = cnt[25] ? _GEN_6276 : _GEN_6139; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6350 = cnt[25] ? _GEN_6277 : _GEN_6140; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6351 = cnt[25] ? _GEN_6278 : _GEN_6141; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6352 = cnt[25] ? _GEN_6279 : _GEN_6142; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6353 = cnt[25] ? _GEN_6280 : _GEN_6143; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6354 = cnt[25] ? _GEN_6281 : _GEN_6144; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6355 = cnt[25] ? _GEN_6282 : _GEN_6145; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6356 = cnt[25] ? _GEN_6283 : _GEN_6146; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6357 = cnt[25] ? _GEN_6284 : _GEN_6147; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6358 = cnt[25] ? _GEN_6285 : _GEN_6148; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6359 = cnt[25] ? _GEN_6286 : _GEN_6149; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6360 = cnt[25] ? _GEN_6287 : _GEN_6150; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6361 = cnt[25] ? _GEN_6288 : _GEN_6151; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6362 = cnt[25] ? _GEN_6289 : _GEN_6152; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6363 = cnt[25] ? _GEN_6290 : _GEN_6153; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6364 = cnt[25] ? _GEN_6291 : _GEN_6154; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6365 = cnt[25] ? _GEN_6292 : _GEN_6155; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6366 = cnt[25] ? _GEN_6293 : _GEN_6156; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6367 = cnt[25] ? _GEN_6294 : _GEN_6157; // @[NulCtrlMP.scala 843:29]
  wire [8:0] _T_510 = pgbuf_cpu_pos[11:3] + 9'h5; // @[NulCtrlMP.scala 843:77]
  wire  _GEN_6368 = _GEN_145 | _GEN_6295; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6369 = _GEN_146 | _GEN_6296; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6370 = _GEN_147 | _GEN_6297; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6371 = _GEN_148 | _GEN_6298; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_6372 = 2'h0 == opidx ? 5'hb : _GEN_6299; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6373 = 2'h1 == opidx ? 5'hb : _GEN_6300; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6374 = 2'h2 == opidx ? 5'hb : _GEN_6301; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6375 = 2'h3 == opidx ? 5'hb : _GEN_6302; // @[NulCtrlMP.scala 352:{28,28}]
  wire [63:0] _GEN_6376 = 6'h0 == _T_510[5:0] ? _GEN_1349 : _GEN_6304; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6377 = 6'h1 == _T_510[5:0] ? _GEN_1349 : _GEN_6305; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6378 = 6'h2 == _T_510[5:0] ? _GEN_1349 : _GEN_6306; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6379 = 6'h3 == _T_510[5:0] ? _GEN_1349 : _GEN_6307; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6380 = 6'h4 == _T_510[5:0] ? _GEN_1349 : _GEN_6308; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6381 = 6'h5 == _T_510[5:0] ? _GEN_1349 : _GEN_6309; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6382 = 6'h6 == _T_510[5:0] ? _GEN_1349 : _GEN_6310; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6383 = 6'h7 == _T_510[5:0] ? _GEN_1349 : _GEN_6311; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6384 = 6'h8 == _T_510[5:0] ? _GEN_1349 : _GEN_6312; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6385 = 6'h9 == _T_510[5:0] ? _GEN_1349 : _GEN_6313; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6386 = 6'ha == _T_510[5:0] ? _GEN_1349 : _GEN_6314; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6387 = 6'hb == _T_510[5:0] ? _GEN_1349 : _GEN_6315; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6388 = 6'hc == _T_510[5:0] ? _GEN_1349 : _GEN_6316; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6389 = 6'hd == _T_510[5:0] ? _GEN_1349 : _GEN_6317; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6390 = 6'he == _T_510[5:0] ? _GEN_1349 : _GEN_6318; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6391 = 6'hf == _T_510[5:0] ? _GEN_1349 : _GEN_6319; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6392 = 6'h10 == _T_510[5:0] ? _GEN_1349 : _GEN_6320; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6393 = 6'h11 == _T_510[5:0] ? _GEN_1349 : _GEN_6321; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6394 = 6'h12 == _T_510[5:0] ? _GEN_1349 : _GEN_6322; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6395 = 6'h13 == _T_510[5:0] ? _GEN_1349 : _GEN_6323; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6396 = 6'h14 == _T_510[5:0] ? _GEN_1349 : _GEN_6324; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6397 = 6'h15 == _T_510[5:0] ? _GEN_1349 : _GEN_6325; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6398 = 6'h16 == _T_510[5:0] ? _GEN_1349 : _GEN_6326; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6399 = 6'h17 == _T_510[5:0] ? _GEN_1349 : _GEN_6327; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6400 = 6'h18 == _T_510[5:0] ? _GEN_1349 : _GEN_6328; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6401 = 6'h19 == _T_510[5:0] ? _GEN_1349 : _GEN_6329; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6402 = 6'h1a == _T_510[5:0] ? _GEN_1349 : _GEN_6330; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6403 = 6'h1b == _T_510[5:0] ? _GEN_1349 : _GEN_6331; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6404 = 6'h1c == _T_510[5:0] ? _GEN_1349 : _GEN_6332; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6405 = 6'h1d == _T_510[5:0] ? _GEN_1349 : _GEN_6333; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6406 = 6'h1e == _T_510[5:0] ? _GEN_1349 : _GEN_6334; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6407 = 6'h1f == _T_510[5:0] ? _GEN_1349 : _GEN_6335; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6408 = 6'h20 == _T_510[5:0] ? _GEN_1349 : _GEN_6336; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6409 = 6'h21 == _T_510[5:0] ? _GEN_1349 : _GEN_6337; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6410 = 6'h22 == _T_510[5:0] ? _GEN_1349 : _GEN_6338; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6411 = 6'h23 == _T_510[5:0] ? _GEN_1349 : _GEN_6339; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6412 = 6'h24 == _T_510[5:0] ? _GEN_1349 : _GEN_6340; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6413 = 6'h25 == _T_510[5:0] ? _GEN_1349 : _GEN_6341; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6414 = 6'h26 == _T_510[5:0] ? _GEN_1349 : _GEN_6342; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6415 = 6'h27 == _T_510[5:0] ? _GEN_1349 : _GEN_6343; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6416 = 6'h28 == _T_510[5:0] ? _GEN_1349 : _GEN_6344; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6417 = 6'h29 == _T_510[5:0] ? _GEN_1349 : _GEN_6345; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6418 = 6'h2a == _T_510[5:0] ? _GEN_1349 : _GEN_6346; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6419 = 6'h2b == _T_510[5:0] ? _GEN_1349 : _GEN_6347; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6420 = 6'h2c == _T_510[5:0] ? _GEN_1349 : _GEN_6348; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6421 = 6'h2d == _T_510[5:0] ? _GEN_1349 : _GEN_6349; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6422 = 6'h2e == _T_510[5:0] ? _GEN_1349 : _GEN_6350; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6423 = 6'h2f == _T_510[5:0] ? _GEN_1349 : _GEN_6351; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6424 = 6'h30 == _T_510[5:0] ? _GEN_1349 : _GEN_6352; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6425 = 6'h31 == _T_510[5:0] ? _GEN_1349 : _GEN_6353; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6426 = 6'h32 == _T_510[5:0] ? _GEN_1349 : _GEN_6354; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6427 = 6'h33 == _T_510[5:0] ? _GEN_1349 : _GEN_6355; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6428 = 6'h34 == _T_510[5:0] ? _GEN_1349 : _GEN_6356; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6429 = 6'h35 == _T_510[5:0] ? _GEN_1349 : _GEN_6357; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6430 = 6'h36 == _T_510[5:0] ? _GEN_1349 : _GEN_6358; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6431 = 6'h37 == _T_510[5:0] ? _GEN_1349 : _GEN_6359; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6432 = 6'h38 == _T_510[5:0] ? _GEN_1349 : _GEN_6360; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6433 = 6'h39 == _T_510[5:0] ? _GEN_1349 : _GEN_6361; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6434 = 6'h3a == _T_510[5:0] ? _GEN_1349 : _GEN_6362; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6435 = 6'h3b == _T_510[5:0] ? _GEN_1349 : _GEN_6363; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6436 = 6'h3c == _T_510[5:0] ? _GEN_1349 : _GEN_6364; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6437 = 6'h3d == _T_510[5:0] ? _GEN_1349 : _GEN_6365; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6438 = 6'h3e == _T_510[5:0] ? _GEN_1349 : _GEN_6366; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6439 = 6'h3f == _T_510[5:0] ? _GEN_1349 : _GEN_6367; // @[NulCtrlMP.scala 355:{17,17}]
  wire [128:0] _GEN_6440 = _T_122 ? _cnt_T : _GEN_6303; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_6441 = _T_122 ? _GEN_6376 : _GEN_6304; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6442 = _T_122 ? _GEN_6377 : _GEN_6305; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6443 = _T_122 ? _GEN_6378 : _GEN_6306; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6444 = _T_122 ? _GEN_6379 : _GEN_6307; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6445 = _T_122 ? _GEN_6380 : _GEN_6308; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6446 = _T_122 ? _GEN_6381 : _GEN_6309; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6447 = _T_122 ? _GEN_6382 : _GEN_6310; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6448 = _T_122 ? _GEN_6383 : _GEN_6311; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6449 = _T_122 ? _GEN_6384 : _GEN_6312; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6450 = _T_122 ? _GEN_6385 : _GEN_6313; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6451 = _T_122 ? _GEN_6386 : _GEN_6314; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6452 = _T_122 ? _GEN_6387 : _GEN_6315; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6453 = _T_122 ? _GEN_6388 : _GEN_6316; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6454 = _T_122 ? _GEN_6389 : _GEN_6317; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6455 = _T_122 ? _GEN_6390 : _GEN_6318; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6456 = _T_122 ? _GEN_6391 : _GEN_6319; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6457 = _T_122 ? _GEN_6392 : _GEN_6320; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6458 = _T_122 ? _GEN_6393 : _GEN_6321; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6459 = _T_122 ? _GEN_6394 : _GEN_6322; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6460 = _T_122 ? _GEN_6395 : _GEN_6323; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6461 = _T_122 ? _GEN_6396 : _GEN_6324; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6462 = _T_122 ? _GEN_6397 : _GEN_6325; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6463 = _T_122 ? _GEN_6398 : _GEN_6326; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6464 = _T_122 ? _GEN_6399 : _GEN_6327; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6465 = _T_122 ? _GEN_6400 : _GEN_6328; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6466 = _T_122 ? _GEN_6401 : _GEN_6329; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6467 = _T_122 ? _GEN_6402 : _GEN_6330; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6468 = _T_122 ? _GEN_6403 : _GEN_6331; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6469 = _T_122 ? _GEN_6404 : _GEN_6332; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6470 = _T_122 ? _GEN_6405 : _GEN_6333; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6471 = _T_122 ? _GEN_6406 : _GEN_6334; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6472 = _T_122 ? _GEN_6407 : _GEN_6335; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6473 = _T_122 ? _GEN_6408 : _GEN_6336; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6474 = _T_122 ? _GEN_6409 : _GEN_6337; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6475 = _T_122 ? _GEN_6410 : _GEN_6338; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6476 = _T_122 ? _GEN_6411 : _GEN_6339; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6477 = _T_122 ? _GEN_6412 : _GEN_6340; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6478 = _T_122 ? _GEN_6413 : _GEN_6341; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6479 = _T_122 ? _GEN_6414 : _GEN_6342; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6480 = _T_122 ? _GEN_6415 : _GEN_6343; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6481 = _T_122 ? _GEN_6416 : _GEN_6344; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6482 = _T_122 ? _GEN_6417 : _GEN_6345; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6483 = _T_122 ? _GEN_6418 : _GEN_6346; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6484 = _T_122 ? _GEN_6419 : _GEN_6347; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6485 = _T_122 ? _GEN_6420 : _GEN_6348; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6486 = _T_122 ? _GEN_6421 : _GEN_6349; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6487 = _T_122 ? _GEN_6422 : _GEN_6350; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6488 = _T_122 ? _GEN_6423 : _GEN_6351; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6489 = _T_122 ? _GEN_6424 : _GEN_6352; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6490 = _T_122 ? _GEN_6425 : _GEN_6353; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6491 = _T_122 ? _GEN_6426 : _GEN_6354; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6492 = _T_122 ? _GEN_6427 : _GEN_6355; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6493 = _T_122 ? _GEN_6428 : _GEN_6356; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6494 = _T_122 ? _GEN_6429 : _GEN_6357; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6495 = _T_122 ? _GEN_6430 : _GEN_6358; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6496 = _T_122 ? _GEN_6431 : _GEN_6359; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6497 = _T_122 ? _GEN_6432 : _GEN_6360; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6498 = _T_122 ? _GEN_6433 : _GEN_6361; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6499 = _T_122 ? _GEN_6434 : _GEN_6362; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6500 = _T_122 ? _GEN_6435 : _GEN_6363; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6501 = _T_122 ? _GEN_6436 : _GEN_6364; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6502 = _T_122 ? _GEN_6437 : _GEN_6365; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6503 = _T_122 ? _GEN_6438 : _GEN_6366; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6504 = _T_122 ? _GEN_6439 : _GEN_6367; // @[NulCtrlMP.scala 353:36]
  wire  _GEN_6505 = cnt[26] ? _GEN_6368 : _GEN_6295; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6506 = cnt[26] ? _GEN_6369 : _GEN_6296; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6507 = cnt[26] ? _GEN_6370 : _GEN_6297; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6508 = cnt[26] ? _GEN_6371 : _GEN_6298; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6509 = cnt[26] ? _GEN_6372 : _GEN_6299; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6510 = cnt[26] ? _GEN_6373 : _GEN_6300; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6511 = cnt[26] ? _GEN_6374 : _GEN_6301; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6512 = cnt[26] ? _GEN_6375 : _GEN_6302; // @[NulCtrlMP.scala 843:29]
  wire [128:0] _GEN_6513 = cnt[26] ? _GEN_6440 : _GEN_6303; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6514 = cnt[26] ? _GEN_6441 : _GEN_6304; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6515 = cnt[26] ? _GEN_6442 : _GEN_6305; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6516 = cnt[26] ? _GEN_6443 : _GEN_6306; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6517 = cnt[26] ? _GEN_6444 : _GEN_6307; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6518 = cnt[26] ? _GEN_6445 : _GEN_6308; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6519 = cnt[26] ? _GEN_6446 : _GEN_6309; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6520 = cnt[26] ? _GEN_6447 : _GEN_6310; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6521 = cnt[26] ? _GEN_6448 : _GEN_6311; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6522 = cnt[26] ? _GEN_6449 : _GEN_6312; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6523 = cnt[26] ? _GEN_6450 : _GEN_6313; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6524 = cnt[26] ? _GEN_6451 : _GEN_6314; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6525 = cnt[26] ? _GEN_6452 : _GEN_6315; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6526 = cnt[26] ? _GEN_6453 : _GEN_6316; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6527 = cnt[26] ? _GEN_6454 : _GEN_6317; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6528 = cnt[26] ? _GEN_6455 : _GEN_6318; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6529 = cnt[26] ? _GEN_6456 : _GEN_6319; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6530 = cnt[26] ? _GEN_6457 : _GEN_6320; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6531 = cnt[26] ? _GEN_6458 : _GEN_6321; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6532 = cnt[26] ? _GEN_6459 : _GEN_6322; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6533 = cnt[26] ? _GEN_6460 : _GEN_6323; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6534 = cnt[26] ? _GEN_6461 : _GEN_6324; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6535 = cnt[26] ? _GEN_6462 : _GEN_6325; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6536 = cnt[26] ? _GEN_6463 : _GEN_6326; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6537 = cnt[26] ? _GEN_6464 : _GEN_6327; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6538 = cnt[26] ? _GEN_6465 : _GEN_6328; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6539 = cnt[26] ? _GEN_6466 : _GEN_6329; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6540 = cnt[26] ? _GEN_6467 : _GEN_6330; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6541 = cnt[26] ? _GEN_6468 : _GEN_6331; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6542 = cnt[26] ? _GEN_6469 : _GEN_6332; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6543 = cnt[26] ? _GEN_6470 : _GEN_6333; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6544 = cnt[26] ? _GEN_6471 : _GEN_6334; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6545 = cnt[26] ? _GEN_6472 : _GEN_6335; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6546 = cnt[26] ? _GEN_6473 : _GEN_6336; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6547 = cnt[26] ? _GEN_6474 : _GEN_6337; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6548 = cnt[26] ? _GEN_6475 : _GEN_6338; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6549 = cnt[26] ? _GEN_6476 : _GEN_6339; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6550 = cnt[26] ? _GEN_6477 : _GEN_6340; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6551 = cnt[26] ? _GEN_6478 : _GEN_6341; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6552 = cnt[26] ? _GEN_6479 : _GEN_6342; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6553 = cnt[26] ? _GEN_6480 : _GEN_6343; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6554 = cnt[26] ? _GEN_6481 : _GEN_6344; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6555 = cnt[26] ? _GEN_6482 : _GEN_6345; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6556 = cnt[26] ? _GEN_6483 : _GEN_6346; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6557 = cnt[26] ? _GEN_6484 : _GEN_6347; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6558 = cnt[26] ? _GEN_6485 : _GEN_6348; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6559 = cnt[26] ? _GEN_6486 : _GEN_6349; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6560 = cnt[26] ? _GEN_6487 : _GEN_6350; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6561 = cnt[26] ? _GEN_6488 : _GEN_6351; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6562 = cnt[26] ? _GEN_6489 : _GEN_6352; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6563 = cnt[26] ? _GEN_6490 : _GEN_6353; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6564 = cnt[26] ? _GEN_6491 : _GEN_6354; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6565 = cnt[26] ? _GEN_6492 : _GEN_6355; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6566 = cnt[26] ? _GEN_6493 : _GEN_6356; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6567 = cnt[26] ? _GEN_6494 : _GEN_6357; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6568 = cnt[26] ? _GEN_6495 : _GEN_6358; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6569 = cnt[26] ? _GEN_6496 : _GEN_6359; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6570 = cnt[26] ? _GEN_6497 : _GEN_6360; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6571 = cnt[26] ? _GEN_6498 : _GEN_6361; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6572 = cnt[26] ? _GEN_6499 : _GEN_6362; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6573 = cnt[26] ? _GEN_6500 : _GEN_6363; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6574 = cnt[26] ? _GEN_6501 : _GEN_6364; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6575 = cnt[26] ? _GEN_6502 : _GEN_6365; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6576 = cnt[26] ? _GEN_6503 : _GEN_6366; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6577 = cnt[26] ? _GEN_6504 : _GEN_6367; // @[NulCtrlMP.scala 843:29]
  wire [8:0] _T_516 = pgbuf_cpu_pos[11:3] + 9'h6; // @[NulCtrlMP.scala 843:77]
  wire  _GEN_6578 = _GEN_145 | _GEN_6505; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6579 = _GEN_146 | _GEN_6506; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6580 = _GEN_147 | _GEN_6507; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6581 = _GEN_148 | _GEN_6508; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_6582 = 2'h0 == opidx ? 5'hc : _GEN_6509; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6583 = 2'h1 == opidx ? 5'hc : _GEN_6510; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6584 = 2'h2 == opidx ? 5'hc : _GEN_6511; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6585 = 2'h3 == opidx ? 5'hc : _GEN_6512; // @[NulCtrlMP.scala 352:{28,28}]
  wire [63:0] _GEN_6586 = 6'h0 == _T_516[5:0] ? _GEN_1349 : _GEN_6514; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6587 = 6'h1 == _T_516[5:0] ? _GEN_1349 : _GEN_6515; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6588 = 6'h2 == _T_516[5:0] ? _GEN_1349 : _GEN_6516; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6589 = 6'h3 == _T_516[5:0] ? _GEN_1349 : _GEN_6517; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6590 = 6'h4 == _T_516[5:0] ? _GEN_1349 : _GEN_6518; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6591 = 6'h5 == _T_516[5:0] ? _GEN_1349 : _GEN_6519; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6592 = 6'h6 == _T_516[5:0] ? _GEN_1349 : _GEN_6520; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6593 = 6'h7 == _T_516[5:0] ? _GEN_1349 : _GEN_6521; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6594 = 6'h8 == _T_516[5:0] ? _GEN_1349 : _GEN_6522; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6595 = 6'h9 == _T_516[5:0] ? _GEN_1349 : _GEN_6523; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6596 = 6'ha == _T_516[5:0] ? _GEN_1349 : _GEN_6524; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6597 = 6'hb == _T_516[5:0] ? _GEN_1349 : _GEN_6525; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6598 = 6'hc == _T_516[5:0] ? _GEN_1349 : _GEN_6526; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6599 = 6'hd == _T_516[5:0] ? _GEN_1349 : _GEN_6527; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6600 = 6'he == _T_516[5:0] ? _GEN_1349 : _GEN_6528; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6601 = 6'hf == _T_516[5:0] ? _GEN_1349 : _GEN_6529; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6602 = 6'h10 == _T_516[5:0] ? _GEN_1349 : _GEN_6530; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6603 = 6'h11 == _T_516[5:0] ? _GEN_1349 : _GEN_6531; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6604 = 6'h12 == _T_516[5:0] ? _GEN_1349 : _GEN_6532; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6605 = 6'h13 == _T_516[5:0] ? _GEN_1349 : _GEN_6533; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6606 = 6'h14 == _T_516[5:0] ? _GEN_1349 : _GEN_6534; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6607 = 6'h15 == _T_516[5:0] ? _GEN_1349 : _GEN_6535; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6608 = 6'h16 == _T_516[5:0] ? _GEN_1349 : _GEN_6536; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6609 = 6'h17 == _T_516[5:0] ? _GEN_1349 : _GEN_6537; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6610 = 6'h18 == _T_516[5:0] ? _GEN_1349 : _GEN_6538; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6611 = 6'h19 == _T_516[5:0] ? _GEN_1349 : _GEN_6539; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6612 = 6'h1a == _T_516[5:0] ? _GEN_1349 : _GEN_6540; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6613 = 6'h1b == _T_516[5:0] ? _GEN_1349 : _GEN_6541; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6614 = 6'h1c == _T_516[5:0] ? _GEN_1349 : _GEN_6542; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6615 = 6'h1d == _T_516[5:0] ? _GEN_1349 : _GEN_6543; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6616 = 6'h1e == _T_516[5:0] ? _GEN_1349 : _GEN_6544; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6617 = 6'h1f == _T_516[5:0] ? _GEN_1349 : _GEN_6545; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6618 = 6'h20 == _T_516[5:0] ? _GEN_1349 : _GEN_6546; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6619 = 6'h21 == _T_516[5:0] ? _GEN_1349 : _GEN_6547; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6620 = 6'h22 == _T_516[5:0] ? _GEN_1349 : _GEN_6548; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6621 = 6'h23 == _T_516[5:0] ? _GEN_1349 : _GEN_6549; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6622 = 6'h24 == _T_516[5:0] ? _GEN_1349 : _GEN_6550; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6623 = 6'h25 == _T_516[5:0] ? _GEN_1349 : _GEN_6551; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6624 = 6'h26 == _T_516[5:0] ? _GEN_1349 : _GEN_6552; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6625 = 6'h27 == _T_516[5:0] ? _GEN_1349 : _GEN_6553; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6626 = 6'h28 == _T_516[5:0] ? _GEN_1349 : _GEN_6554; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6627 = 6'h29 == _T_516[5:0] ? _GEN_1349 : _GEN_6555; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6628 = 6'h2a == _T_516[5:0] ? _GEN_1349 : _GEN_6556; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6629 = 6'h2b == _T_516[5:0] ? _GEN_1349 : _GEN_6557; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6630 = 6'h2c == _T_516[5:0] ? _GEN_1349 : _GEN_6558; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6631 = 6'h2d == _T_516[5:0] ? _GEN_1349 : _GEN_6559; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6632 = 6'h2e == _T_516[5:0] ? _GEN_1349 : _GEN_6560; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6633 = 6'h2f == _T_516[5:0] ? _GEN_1349 : _GEN_6561; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6634 = 6'h30 == _T_516[5:0] ? _GEN_1349 : _GEN_6562; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6635 = 6'h31 == _T_516[5:0] ? _GEN_1349 : _GEN_6563; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6636 = 6'h32 == _T_516[5:0] ? _GEN_1349 : _GEN_6564; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6637 = 6'h33 == _T_516[5:0] ? _GEN_1349 : _GEN_6565; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6638 = 6'h34 == _T_516[5:0] ? _GEN_1349 : _GEN_6566; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6639 = 6'h35 == _T_516[5:0] ? _GEN_1349 : _GEN_6567; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6640 = 6'h36 == _T_516[5:0] ? _GEN_1349 : _GEN_6568; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6641 = 6'h37 == _T_516[5:0] ? _GEN_1349 : _GEN_6569; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6642 = 6'h38 == _T_516[5:0] ? _GEN_1349 : _GEN_6570; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6643 = 6'h39 == _T_516[5:0] ? _GEN_1349 : _GEN_6571; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6644 = 6'h3a == _T_516[5:0] ? _GEN_1349 : _GEN_6572; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6645 = 6'h3b == _T_516[5:0] ? _GEN_1349 : _GEN_6573; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6646 = 6'h3c == _T_516[5:0] ? _GEN_1349 : _GEN_6574; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6647 = 6'h3d == _T_516[5:0] ? _GEN_1349 : _GEN_6575; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6648 = 6'h3e == _T_516[5:0] ? _GEN_1349 : _GEN_6576; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6649 = 6'h3f == _T_516[5:0] ? _GEN_1349 : _GEN_6577; // @[NulCtrlMP.scala 355:{17,17}]
  wire [128:0] _GEN_6650 = _T_122 ? _cnt_T : _GEN_6513; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_6651 = _T_122 ? _GEN_6586 : _GEN_6514; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6652 = _T_122 ? _GEN_6587 : _GEN_6515; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6653 = _T_122 ? _GEN_6588 : _GEN_6516; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6654 = _T_122 ? _GEN_6589 : _GEN_6517; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6655 = _T_122 ? _GEN_6590 : _GEN_6518; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6656 = _T_122 ? _GEN_6591 : _GEN_6519; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6657 = _T_122 ? _GEN_6592 : _GEN_6520; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6658 = _T_122 ? _GEN_6593 : _GEN_6521; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6659 = _T_122 ? _GEN_6594 : _GEN_6522; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6660 = _T_122 ? _GEN_6595 : _GEN_6523; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6661 = _T_122 ? _GEN_6596 : _GEN_6524; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6662 = _T_122 ? _GEN_6597 : _GEN_6525; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6663 = _T_122 ? _GEN_6598 : _GEN_6526; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6664 = _T_122 ? _GEN_6599 : _GEN_6527; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6665 = _T_122 ? _GEN_6600 : _GEN_6528; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6666 = _T_122 ? _GEN_6601 : _GEN_6529; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6667 = _T_122 ? _GEN_6602 : _GEN_6530; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6668 = _T_122 ? _GEN_6603 : _GEN_6531; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6669 = _T_122 ? _GEN_6604 : _GEN_6532; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6670 = _T_122 ? _GEN_6605 : _GEN_6533; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6671 = _T_122 ? _GEN_6606 : _GEN_6534; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6672 = _T_122 ? _GEN_6607 : _GEN_6535; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6673 = _T_122 ? _GEN_6608 : _GEN_6536; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6674 = _T_122 ? _GEN_6609 : _GEN_6537; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6675 = _T_122 ? _GEN_6610 : _GEN_6538; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6676 = _T_122 ? _GEN_6611 : _GEN_6539; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6677 = _T_122 ? _GEN_6612 : _GEN_6540; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6678 = _T_122 ? _GEN_6613 : _GEN_6541; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6679 = _T_122 ? _GEN_6614 : _GEN_6542; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6680 = _T_122 ? _GEN_6615 : _GEN_6543; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6681 = _T_122 ? _GEN_6616 : _GEN_6544; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6682 = _T_122 ? _GEN_6617 : _GEN_6545; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6683 = _T_122 ? _GEN_6618 : _GEN_6546; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6684 = _T_122 ? _GEN_6619 : _GEN_6547; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6685 = _T_122 ? _GEN_6620 : _GEN_6548; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6686 = _T_122 ? _GEN_6621 : _GEN_6549; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6687 = _T_122 ? _GEN_6622 : _GEN_6550; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6688 = _T_122 ? _GEN_6623 : _GEN_6551; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6689 = _T_122 ? _GEN_6624 : _GEN_6552; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6690 = _T_122 ? _GEN_6625 : _GEN_6553; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6691 = _T_122 ? _GEN_6626 : _GEN_6554; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6692 = _T_122 ? _GEN_6627 : _GEN_6555; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6693 = _T_122 ? _GEN_6628 : _GEN_6556; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6694 = _T_122 ? _GEN_6629 : _GEN_6557; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6695 = _T_122 ? _GEN_6630 : _GEN_6558; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6696 = _T_122 ? _GEN_6631 : _GEN_6559; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6697 = _T_122 ? _GEN_6632 : _GEN_6560; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6698 = _T_122 ? _GEN_6633 : _GEN_6561; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6699 = _T_122 ? _GEN_6634 : _GEN_6562; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6700 = _T_122 ? _GEN_6635 : _GEN_6563; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6701 = _T_122 ? _GEN_6636 : _GEN_6564; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6702 = _T_122 ? _GEN_6637 : _GEN_6565; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6703 = _T_122 ? _GEN_6638 : _GEN_6566; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6704 = _T_122 ? _GEN_6639 : _GEN_6567; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6705 = _T_122 ? _GEN_6640 : _GEN_6568; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6706 = _T_122 ? _GEN_6641 : _GEN_6569; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6707 = _T_122 ? _GEN_6642 : _GEN_6570; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6708 = _T_122 ? _GEN_6643 : _GEN_6571; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6709 = _T_122 ? _GEN_6644 : _GEN_6572; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6710 = _T_122 ? _GEN_6645 : _GEN_6573; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6711 = _T_122 ? _GEN_6646 : _GEN_6574; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6712 = _T_122 ? _GEN_6647 : _GEN_6575; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6713 = _T_122 ? _GEN_6648 : _GEN_6576; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6714 = _T_122 ? _GEN_6649 : _GEN_6577; // @[NulCtrlMP.scala 353:36]
  wire  _GEN_6715 = cnt[27] ? _GEN_6578 : _GEN_6505; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6716 = cnt[27] ? _GEN_6579 : _GEN_6506; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6717 = cnt[27] ? _GEN_6580 : _GEN_6507; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6718 = cnt[27] ? _GEN_6581 : _GEN_6508; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6719 = cnt[27] ? _GEN_6582 : _GEN_6509; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6720 = cnt[27] ? _GEN_6583 : _GEN_6510; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6721 = cnt[27] ? _GEN_6584 : _GEN_6511; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6722 = cnt[27] ? _GEN_6585 : _GEN_6512; // @[NulCtrlMP.scala 843:29]
  wire [128:0] _GEN_6723 = cnt[27] ? _GEN_6650 : _GEN_6513; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6724 = cnt[27] ? _GEN_6651 : _GEN_6514; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6725 = cnt[27] ? _GEN_6652 : _GEN_6515; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6726 = cnt[27] ? _GEN_6653 : _GEN_6516; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6727 = cnt[27] ? _GEN_6654 : _GEN_6517; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6728 = cnt[27] ? _GEN_6655 : _GEN_6518; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6729 = cnt[27] ? _GEN_6656 : _GEN_6519; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6730 = cnt[27] ? _GEN_6657 : _GEN_6520; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6731 = cnt[27] ? _GEN_6658 : _GEN_6521; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6732 = cnt[27] ? _GEN_6659 : _GEN_6522; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6733 = cnt[27] ? _GEN_6660 : _GEN_6523; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6734 = cnt[27] ? _GEN_6661 : _GEN_6524; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6735 = cnt[27] ? _GEN_6662 : _GEN_6525; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6736 = cnt[27] ? _GEN_6663 : _GEN_6526; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6737 = cnt[27] ? _GEN_6664 : _GEN_6527; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6738 = cnt[27] ? _GEN_6665 : _GEN_6528; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6739 = cnt[27] ? _GEN_6666 : _GEN_6529; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6740 = cnt[27] ? _GEN_6667 : _GEN_6530; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6741 = cnt[27] ? _GEN_6668 : _GEN_6531; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6742 = cnt[27] ? _GEN_6669 : _GEN_6532; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6743 = cnt[27] ? _GEN_6670 : _GEN_6533; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6744 = cnt[27] ? _GEN_6671 : _GEN_6534; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6745 = cnt[27] ? _GEN_6672 : _GEN_6535; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6746 = cnt[27] ? _GEN_6673 : _GEN_6536; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6747 = cnt[27] ? _GEN_6674 : _GEN_6537; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6748 = cnt[27] ? _GEN_6675 : _GEN_6538; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6749 = cnt[27] ? _GEN_6676 : _GEN_6539; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6750 = cnt[27] ? _GEN_6677 : _GEN_6540; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6751 = cnt[27] ? _GEN_6678 : _GEN_6541; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6752 = cnt[27] ? _GEN_6679 : _GEN_6542; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6753 = cnt[27] ? _GEN_6680 : _GEN_6543; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6754 = cnt[27] ? _GEN_6681 : _GEN_6544; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6755 = cnt[27] ? _GEN_6682 : _GEN_6545; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6756 = cnt[27] ? _GEN_6683 : _GEN_6546; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6757 = cnt[27] ? _GEN_6684 : _GEN_6547; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6758 = cnt[27] ? _GEN_6685 : _GEN_6548; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6759 = cnt[27] ? _GEN_6686 : _GEN_6549; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6760 = cnt[27] ? _GEN_6687 : _GEN_6550; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6761 = cnt[27] ? _GEN_6688 : _GEN_6551; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6762 = cnt[27] ? _GEN_6689 : _GEN_6552; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6763 = cnt[27] ? _GEN_6690 : _GEN_6553; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6764 = cnt[27] ? _GEN_6691 : _GEN_6554; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6765 = cnt[27] ? _GEN_6692 : _GEN_6555; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6766 = cnt[27] ? _GEN_6693 : _GEN_6556; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6767 = cnt[27] ? _GEN_6694 : _GEN_6557; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6768 = cnt[27] ? _GEN_6695 : _GEN_6558; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6769 = cnt[27] ? _GEN_6696 : _GEN_6559; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6770 = cnt[27] ? _GEN_6697 : _GEN_6560; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6771 = cnt[27] ? _GEN_6698 : _GEN_6561; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6772 = cnt[27] ? _GEN_6699 : _GEN_6562; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6773 = cnt[27] ? _GEN_6700 : _GEN_6563; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6774 = cnt[27] ? _GEN_6701 : _GEN_6564; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6775 = cnt[27] ? _GEN_6702 : _GEN_6565; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6776 = cnt[27] ? _GEN_6703 : _GEN_6566; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6777 = cnt[27] ? _GEN_6704 : _GEN_6567; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6778 = cnt[27] ? _GEN_6705 : _GEN_6568; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6779 = cnt[27] ? _GEN_6706 : _GEN_6569; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6780 = cnt[27] ? _GEN_6707 : _GEN_6570; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6781 = cnt[27] ? _GEN_6708 : _GEN_6571; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6782 = cnt[27] ? _GEN_6709 : _GEN_6572; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6783 = cnt[27] ? _GEN_6710 : _GEN_6573; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6784 = cnt[27] ? _GEN_6711 : _GEN_6574; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6785 = cnt[27] ? _GEN_6712 : _GEN_6575; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6786 = cnt[27] ? _GEN_6713 : _GEN_6576; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6787 = cnt[27] ? _GEN_6714 : _GEN_6577; // @[NulCtrlMP.scala 843:29]
  wire [8:0] _T_522 = pgbuf_cpu_pos[11:3] + 9'h7; // @[NulCtrlMP.scala 843:77]
  wire  _GEN_6788 = _GEN_145 | _GEN_6715; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6789 = _GEN_146 | _GEN_6716; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6790 = _GEN_147 | _GEN_6717; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_6791 = _GEN_148 | _GEN_6718; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_6792 = 2'h0 == opidx ? 5'hd : _GEN_6719; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6793 = 2'h1 == opidx ? 5'hd : _GEN_6720; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6794 = 2'h2 == opidx ? 5'hd : _GEN_6721; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_6795 = 2'h3 == opidx ? 5'hd : _GEN_6722; // @[NulCtrlMP.scala 352:{28,28}]
  wire [63:0] _GEN_6796 = 6'h0 == _T_522[5:0] ? _GEN_1349 : _GEN_6724; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6797 = 6'h1 == _T_522[5:0] ? _GEN_1349 : _GEN_6725; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6798 = 6'h2 == _T_522[5:0] ? _GEN_1349 : _GEN_6726; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6799 = 6'h3 == _T_522[5:0] ? _GEN_1349 : _GEN_6727; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6800 = 6'h4 == _T_522[5:0] ? _GEN_1349 : _GEN_6728; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6801 = 6'h5 == _T_522[5:0] ? _GEN_1349 : _GEN_6729; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6802 = 6'h6 == _T_522[5:0] ? _GEN_1349 : _GEN_6730; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6803 = 6'h7 == _T_522[5:0] ? _GEN_1349 : _GEN_6731; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6804 = 6'h8 == _T_522[5:0] ? _GEN_1349 : _GEN_6732; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6805 = 6'h9 == _T_522[5:0] ? _GEN_1349 : _GEN_6733; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6806 = 6'ha == _T_522[5:0] ? _GEN_1349 : _GEN_6734; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6807 = 6'hb == _T_522[5:0] ? _GEN_1349 : _GEN_6735; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6808 = 6'hc == _T_522[5:0] ? _GEN_1349 : _GEN_6736; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6809 = 6'hd == _T_522[5:0] ? _GEN_1349 : _GEN_6737; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6810 = 6'he == _T_522[5:0] ? _GEN_1349 : _GEN_6738; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6811 = 6'hf == _T_522[5:0] ? _GEN_1349 : _GEN_6739; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6812 = 6'h10 == _T_522[5:0] ? _GEN_1349 : _GEN_6740; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6813 = 6'h11 == _T_522[5:0] ? _GEN_1349 : _GEN_6741; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6814 = 6'h12 == _T_522[5:0] ? _GEN_1349 : _GEN_6742; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6815 = 6'h13 == _T_522[5:0] ? _GEN_1349 : _GEN_6743; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6816 = 6'h14 == _T_522[5:0] ? _GEN_1349 : _GEN_6744; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6817 = 6'h15 == _T_522[5:0] ? _GEN_1349 : _GEN_6745; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6818 = 6'h16 == _T_522[5:0] ? _GEN_1349 : _GEN_6746; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6819 = 6'h17 == _T_522[5:0] ? _GEN_1349 : _GEN_6747; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6820 = 6'h18 == _T_522[5:0] ? _GEN_1349 : _GEN_6748; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6821 = 6'h19 == _T_522[5:0] ? _GEN_1349 : _GEN_6749; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6822 = 6'h1a == _T_522[5:0] ? _GEN_1349 : _GEN_6750; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6823 = 6'h1b == _T_522[5:0] ? _GEN_1349 : _GEN_6751; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6824 = 6'h1c == _T_522[5:0] ? _GEN_1349 : _GEN_6752; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6825 = 6'h1d == _T_522[5:0] ? _GEN_1349 : _GEN_6753; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6826 = 6'h1e == _T_522[5:0] ? _GEN_1349 : _GEN_6754; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6827 = 6'h1f == _T_522[5:0] ? _GEN_1349 : _GEN_6755; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6828 = 6'h20 == _T_522[5:0] ? _GEN_1349 : _GEN_6756; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6829 = 6'h21 == _T_522[5:0] ? _GEN_1349 : _GEN_6757; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6830 = 6'h22 == _T_522[5:0] ? _GEN_1349 : _GEN_6758; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6831 = 6'h23 == _T_522[5:0] ? _GEN_1349 : _GEN_6759; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6832 = 6'h24 == _T_522[5:0] ? _GEN_1349 : _GEN_6760; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6833 = 6'h25 == _T_522[5:0] ? _GEN_1349 : _GEN_6761; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6834 = 6'h26 == _T_522[5:0] ? _GEN_1349 : _GEN_6762; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6835 = 6'h27 == _T_522[5:0] ? _GEN_1349 : _GEN_6763; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6836 = 6'h28 == _T_522[5:0] ? _GEN_1349 : _GEN_6764; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6837 = 6'h29 == _T_522[5:0] ? _GEN_1349 : _GEN_6765; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6838 = 6'h2a == _T_522[5:0] ? _GEN_1349 : _GEN_6766; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6839 = 6'h2b == _T_522[5:0] ? _GEN_1349 : _GEN_6767; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6840 = 6'h2c == _T_522[5:0] ? _GEN_1349 : _GEN_6768; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6841 = 6'h2d == _T_522[5:0] ? _GEN_1349 : _GEN_6769; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6842 = 6'h2e == _T_522[5:0] ? _GEN_1349 : _GEN_6770; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6843 = 6'h2f == _T_522[5:0] ? _GEN_1349 : _GEN_6771; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6844 = 6'h30 == _T_522[5:0] ? _GEN_1349 : _GEN_6772; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6845 = 6'h31 == _T_522[5:0] ? _GEN_1349 : _GEN_6773; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6846 = 6'h32 == _T_522[5:0] ? _GEN_1349 : _GEN_6774; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6847 = 6'h33 == _T_522[5:0] ? _GEN_1349 : _GEN_6775; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6848 = 6'h34 == _T_522[5:0] ? _GEN_1349 : _GEN_6776; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6849 = 6'h35 == _T_522[5:0] ? _GEN_1349 : _GEN_6777; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6850 = 6'h36 == _T_522[5:0] ? _GEN_1349 : _GEN_6778; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6851 = 6'h37 == _T_522[5:0] ? _GEN_1349 : _GEN_6779; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6852 = 6'h38 == _T_522[5:0] ? _GEN_1349 : _GEN_6780; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6853 = 6'h39 == _T_522[5:0] ? _GEN_1349 : _GEN_6781; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6854 = 6'h3a == _T_522[5:0] ? _GEN_1349 : _GEN_6782; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6855 = 6'h3b == _T_522[5:0] ? _GEN_1349 : _GEN_6783; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6856 = 6'h3c == _T_522[5:0] ? _GEN_1349 : _GEN_6784; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6857 = 6'h3d == _T_522[5:0] ? _GEN_1349 : _GEN_6785; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6858 = 6'h3e == _T_522[5:0] ? _GEN_1349 : _GEN_6786; // @[NulCtrlMP.scala 355:{17,17}]
  wire [63:0] _GEN_6859 = 6'h3f == _T_522[5:0] ? _GEN_1349 : _GEN_6787; // @[NulCtrlMP.scala 355:{17,17}]
  wire [128:0] _GEN_6860 = _T_122 ? _cnt_T : _GEN_6723; // @[NulCtrlMP.scala 353:36 354:17]
  wire [63:0] _GEN_6861 = _T_122 ? _GEN_6796 : _GEN_6724; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6862 = _T_122 ? _GEN_6797 : _GEN_6725; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6863 = _T_122 ? _GEN_6798 : _GEN_6726; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6864 = _T_122 ? _GEN_6799 : _GEN_6727; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6865 = _T_122 ? _GEN_6800 : _GEN_6728; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6866 = _T_122 ? _GEN_6801 : _GEN_6729; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6867 = _T_122 ? _GEN_6802 : _GEN_6730; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6868 = _T_122 ? _GEN_6803 : _GEN_6731; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6869 = _T_122 ? _GEN_6804 : _GEN_6732; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6870 = _T_122 ? _GEN_6805 : _GEN_6733; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6871 = _T_122 ? _GEN_6806 : _GEN_6734; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6872 = _T_122 ? _GEN_6807 : _GEN_6735; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6873 = _T_122 ? _GEN_6808 : _GEN_6736; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6874 = _T_122 ? _GEN_6809 : _GEN_6737; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6875 = _T_122 ? _GEN_6810 : _GEN_6738; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6876 = _T_122 ? _GEN_6811 : _GEN_6739; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6877 = _T_122 ? _GEN_6812 : _GEN_6740; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6878 = _T_122 ? _GEN_6813 : _GEN_6741; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6879 = _T_122 ? _GEN_6814 : _GEN_6742; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6880 = _T_122 ? _GEN_6815 : _GEN_6743; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6881 = _T_122 ? _GEN_6816 : _GEN_6744; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6882 = _T_122 ? _GEN_6817 : _GEN_6745; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6883 = _T_122 ? _GEN_6818 : _GEN_6746; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6884 = _T_122 ? _GEN_6819 : _GEN_6747; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6885 = _T_122 ? _GEN_6820 : _GEN_6748; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6886 = _T_122 ? _GEN_6821 : _GEN_6749; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6887 = _T_122 ? _GEN_6822 : _GEN_6750; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6888 = _T_122 ? _GEN_6823 : _GEN_6751; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6889 = _T_122 ? _GEN_6824 : _GEN_6752; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6890 = _T_122 ? _GEN_6825 : _GEN_6753; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6891 = _T_122 ? _GEN_6826 : _GEN_6754; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6892 = _T_122 ? _GEN_6827 : _GEN_6755; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6893 = _T_122 ? _GEN_6828 : _GEN_6756; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6894 = _T_122 ? _GEN_6829 : _GEN_6757; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6895 = _T_122 ? _GEN_6830 : _GEN_6758; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6896 = _T_122 ? _GEN_6831 : _GEN_6759; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6897 = _T_122 ? _GEN_6832 : _GEN_6760; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6898 = _T_122 ? _GEN_6833 : _GEN_6761; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6899 = _T_122 ? _GEN_6834 : _GEN_6762; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6900 = _T_122 ? _GEN_6835 : _GEN_6763; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6901 = _T_122 ? _GEN_6836 : _GEN_6764; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6902 = _T_122 ? _GEN_6837 : _GEN_6765; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6903 = _T_122 ? _GEN_6838 : _GEN_6766; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6904 = _T_122 ? _GEN_6839 : _GEN_6767; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6905 = _T_122 ? _GEN_6840 : _GEN_6768; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6906 = _T_122 ? _GEN_6841 : _GEN_6769; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6907 = _T_122 ? _GEN_6842 : _GEN_6770; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6908 = _T_122 ? _GEN_6843 : _GEN_6771; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6909 = _T_122 ? _GEN_6844 : _GEN_6772; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6910 = _T_122 ? _GEN_6845 : _GEN_6773; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6911 = _T_122 ? _GEN_6846 : _GEN_6774; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6912 = _T_122 ? _GEN_6847 : _GEN_6775; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6913 = _T_122 ? _GEN_6848 : _GEN_6776; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6914 = _T_122 ? _GEN_6849 : _GEN_6777; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6915 = _T_122 ? _GEN_6850 : _GEN_6778; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6916 = _T_122 ? _GEN_6851 : _GEN_6779; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6917 = _T_122 ? _GEN_6852 : _GEN_6780; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6918 = _T_122 ? _GEN_6853 : _GEN_6781; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6919 = _T_122 ? _GEN_6854 : _GEN_6782; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6920 = _T_122 ? _GEN_6855 : _GEN_6783; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6921 = _T_122 ? _GEN_6856 : _GEN_6784; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6922 = _T_122 ? _GEN_6857 : _GEN_6785; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6923 = _T_122 ? _GEN_6858 : _GEN_6786; // @[NulCtrlMP.scala 353:36]
  wire [63:0] _GEN_6924 = _T_122 ? _GEN_6859 : _GEN_6787; // @[NulCtrlMP.scala 353:36]
  wire  _GEN_6925 = cnt[28] ? _GEN_6788 : _GEN_6715; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6926 = cnt[28] ? _GEN_6789 : _GEN_6716; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6927 = cnt[28] ? _GEN_6790 : _GEN_6717; // @[NulCtrlMP.scala 843:29]
  wire  _GEN_6928 = cnt[28] ? _GEN_6791 : _GEN_6718; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6929 = cnt[28] ? _GEN_6792 : _GEN_6719; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6930 = cnt[28] ? _GEN_6793 : _GEN_6720; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6931 = cnt[28] ? _GEN_6794 : _GEN_6721; // @[NulCtrlMP.scala 843:29]
  wire [4:0] _GEN_6932 = cnt[28] ? _GEN_6795 : _GEN_6722; // @[NulCtrlMP.scala 843:29]
  wire [128:0] _GEN_6933 = cnt[28] ? _GEN_6860 : _GEN_6723; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6934 = cnt[28] ? _GEN_6861 : _GEN_6724; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6935 = cnt[28] ? _GEN_6862 : _GEN_6725; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6936 = cnt[28] ? _GEN_6863 : _GEN_6726; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6937 = cnt[28] ? _GEN_6864 : _GEN_6727; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6938 = cnt[28] ? _GEN_6865 : _GEN_6728; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6939 = cnt[28] ? _GEN_6866 : _GEN_6729; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6940 = cnt[28] ? _GEN_6867 : _GEN_6730; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6941 = cnt[28] ? _GEN_6868 : _GEN_6731; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6942 = cnt[28] ? _GEN_6869 : _GEN_6732; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6943 = cnt[28] ? _GEN_6870 : _GEN_6733; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6944 = cnt[28] ? _GEN_6871 : _GEN_6734; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6945 = cnt[28] ? _GEN_6872 : _GEN_6735; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6946 = cnt[28] ? _GEN_6873 : _GEN_6736; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6947 = cnt[28] ? _GEN_6874 : _GEN_6737; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6948 = cnt[28] ? _GEN_6875 : _GEN_6738; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6949 = cnt[28] ? _GEN_6876 : _GEN_6739; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6950 = cnt[28] ? _GEN_6877 : _GEN_6740; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6951 = cnt[28] ? _GEN_6878 : _GEN_6741; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6952 = cnt[28] ? _GEN_6879 : _GEN_6742; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6953 = cnt[28] ? _GEN_6880 : _GEN_6743; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6954 = cnt[28] ? _GEN_6881 : _GEN_6744; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6955 = cnt[28] ? _GEN_6882 : _GEN_6745; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6956 = cnt[28] ? _GEN_6883 : _GEN_6746; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6957 = cnt[28] ? _GEN_6884 : _GEN_6747; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6958 = cnt[28] ? _GEN_6885 : _GEN_6748; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6959 = cnt[28] ? _GEN_6886 : _GEN_6749; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6960 = cnt[28] ? _GEN_6887 : _GEN_6750; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6961 = cnt[28] ? _GEN_6888 : _GEN_6751; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6962 = cnt[28] ? _GEN_6889 : _GEN_6752; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6963 = cnt[28] ? _GEN_6890 : _GEN_6753; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6964 = cnt[28] ? _GEN_6891 : _GEN_6754; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6965 = cnt[28] ? _GEN_6892 : _GEN_6755; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6966 = cnt[28] ? _GEN_6893 : _GEN_6756; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6967 = cnt[28] ? _GEN_6894 : _GEN_6757; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6968 = cnt[28] ? _GEN_6895 : _GEN_6758; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6969 = cnt[28] ? _GEN_6896 : _GEN_6759; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6970 = cnt[28] ? _GEN_6897 : _GEN_6760; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6971 = cnt[28] ? _GEN_6898 : _GEN_6761; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6972 = cnt[28] ? _GEN_6899 : _GEN_6762; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6973 = cnt[28] ? _GEN_6900 : _GEN_6763; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6974 = cnt[28] ? _GEN_6901 : _GEN_6764; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6975 = cnt[28] ? _GEN_6902 : _GEN_6765; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6976 = cnt[28] ? _GEN_6903 : _GEN_6766; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6977 = cnt[28] ? _GEN_6904 : _GEN_6767; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6978 = cnt[28] ? _GEN_6905 : _GEN_6768; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6979 = cnt[28] ? _GEN_6906 : _GEN_6769; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6980 = cnt[28] ? _GEN_6907 : _GEN_6770; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6981 = cnt[28] ? _GEN_6908 : _GEN_6771; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6982 = cnt[28] ? _GEN_6909 : _GEN_6772; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6983 = cnt[28] ? _GEN_6910 : _GEN_6773; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6984 = cnt[28] ? _GEN_6911 : _GEN_6774; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6985 = cnt[28] ? _GEN_6912 : _GEN_6775; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6986 = cnt[28] ? _GEN_6913 : _GEN_6776; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6987 = cnt[28] ? _GEN_6914 : _GEN_6777; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6988 = cnt[28] ? _GEN_6915 : _GEN_6778; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6989 = cnt[28] ? _GEN_6916 : _GEN_6779; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6990 = cnt[28] ? _GEN_6917 : _GEN_6780; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6991 = cnt[28] ? _GEN_6918 : _GEN_6781; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6992 = cnt[28] ? _GEN_6919 : _GEN_6782; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6993 = cnt[28] ? _GEN_6920 : _GEN_6783; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6994 = cnt[28] ? _GEN_6921 : _GEN_6784; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6995 = cnt[28] ? _GEN_6922 : _GEN_6785; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6996 = cnt[28] ? _GEN_6923 : _GEN_6786; // @[NulCtrlMP.scala 843:29]
  wire [63:0] _GEN_6997 = cnt[28] ? _GEN_6924 : _GEN_6787; // @[NulCtrlMP.scala 843:29]
  wire  _T_526 = pgbuf_cpu_pos == 12'h1c0; // @[NulCtrlMP.scala 846:32]
  wire [128:0] _GEN_6998 = pgbuf_cpu_pos == 12'h1c0 ? _cnt_T : 129'h800; // @[NulCtrlMP.scala 846:43 847:21 849:21]
  wire [11:0] _pgbuf_cpu_pos_T_1 = pgbuf_cpu_pos + 12'h40; // @[NulCtrlMP.scala 851:44]
  wire [128:0] _GEN_6999 = cnt[29] ? _GEN_6998 : _GEN_6933; // @[NulCtrlMP.scala 845:23]
  wire [11:0] _GEN_7000 = cnt[29] ? _pgbuf_cpu_pos_T_1 : pgbuf_cpu_pos; // @[NulCtrlMP.scala 845:23 851:27 820:32]
  wire  _GEN_7001 = _GEN_145 | _GEN_5299; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_7002 = _GEN_146 | _GEN_5300; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_7003 = _GEN_147 | _GEN_5301; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_7004 = _GEN_148 | _GEN_5302; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_7005 = 2'h0 == opidx ? 32'h330000f : _GEN_5303; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_7006 = 2'h1 == opidx ? 32'h330000f : _GEN_5304; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_7007 = 2'h2 == opidx ? 32'h330000f : _GEN_5305; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_7008 = 2'h3 == opidx ? 32'h330000f : _GEN_5306; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_7009 = _GEN_1180 ? _cnt_T : _GEN_6999; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_7010 = cnt[30] ? _GEN_7001 : _GEN_5299; // @[NulCtrlMP.scala 853:23]
  wire  _GEN_7011 = cnt[30] ? _GEN_7002 : _GEN_5300; // @[NulCtrlMP.scala 853:23]
  wire  _GEN_7012 = cnt[30] ? _GEN_7003 : _GEN_5301; // @[NulCtrlMP.scala 853:23]
  wire  _GEN_7013 = cnt[30] ? _GEN_7004 : _GEN_5302; // @[NulCtrlMP.scala 853:23]
  wire [31:0] _GEN_7014 = cnt[30] ? _GEN_7005 : _GEN_5303; // @[NulCtrlMP.scala 853:23]
  wire [31:0] _GEN_7015 = cnt[30] ? _GEN_7006 : _GEN_5304; // @[NulCtrlMP.scala 853:23]
  wire [31:0] _GEN_7016 = cnt[30] ? _GEN_7007 : _GEN_5305; // @[NulCtrlMP.scala 853:23]
  wire [31:0] _GEN_7017 = cnt[30] ? _GEN_7008 : _GEN_5306; // @[NulCtrlMP.scala 853:23]
  wire [128:0] _GEN_7018 = cnt[30] ? _GEN_7009 : _GEN_6999; // @[NulCtrlMP.scala 853:23]
  wire  _GEN_7019 = _GEN_145 | _GEN_5313; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_7020 = _GEN_146 | _GEN_5314; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_7021 = _GEN_147 | _GEN_5315; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_7022 = _GEN_148 | _GEN_5316; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_7023 = ~_GEN_1252 ? _cnt_T : _GEN_7018; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_7024 = cnt[31] ? _GEN_7019 : _GEN_5313; // @[NulCtrlMP.scala 854:23]
  wire  _GEN_7025 = cnt[31] ? _GEN_7020 : _GEN_5314; // @[NulCtrlMP.scala 854:23]
  wire  _GEN_7026 = cnt[31] ? _GEN_7021 : _GEN_5315; // @[NulCtrlMP.scala 854:23]
  wire  _GEN_7027 = cnt[31] ? _GEN_7022 : _GEN_5316; // @[NulCtrlMP.scala 854:23]
  wire [128:0] _GEN_7028 = cnt[31] ? _GEN_7023 : _GEN_7018; // @[NulCtrlMP.scala 854:23]
  wire  _GEN_7029 = _GEN_145 | _GEN_5133; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7030 = _GEN_146 | _GEN_5134; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7031 = _GEN_147 | _GEN_5135; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7032 = _GEN_148 | _GEN_5136; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7033 = 2'h0 == opidx ? 5'h5 : _GEN_6929; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7034 = 2'h1 == opidx ? 5'h5 : _GEN_6930; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7035 = 2'h2 == opidx ? 5'h5 : _GEN_6931; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7036 = 2'h3 == opidx ? 5'h5 : _GEN_6932; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7037 = 2'h0 == opidx ? regback_0 : _GEN_5141; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7038 = 2'h1 == opidx ? regback_0 : _GEN_5142; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7039 = 2'h2 == opidx ? regback_0 : _GEN_5143; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7040 = 2'h3 == opidx ? regback_0 : _GEN_5144; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7041 = ~_GEN_1128 ? _cnt_T : _GEN_7028; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7042 = cnt[32] ? _GEN_7029 : _GEN_5133; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7043 = cnt[32] ? _GEN_7030 : _GEN_5134; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7044 = cnt[32] ? _GEN_7031 : _GEN_5135; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7045 = cnt[32] ? _GEN_7032 : _GEN_5136; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7046 = cnt[32] ? _GEN_7033 : _GEN_6929; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7047 = cnt[32] ? _GEN_7034 : _GEN_6930; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7048 = cnt[32] ? _GEN_7035 : _GEN_6931; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7049 = cnt[32] ? _GEN_7036 : _GEN_6932; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7050 = cnt[32] ? _GEN_7037 : _GEN_5141; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7051 = cnt[32] ? _GEN_7038 : _GEN_5142; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7052 = cnt[32] ? _GEN_7039 : _GEN_5143; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7053 = cnt[32] ? _GEN_7040 : _GEN_5144; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7054 = cnt[32] ? _GEN_7041 : _GEN_7028; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7055 = _GEN_145 | _GEN_7042; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7056 = _GEN_146 | _GEN_7043; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7057 = _GEN_147 | _GEN_7044; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7058 = _GEN_148 | _GEN_7045; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7059 = 2'h0 == opidx ? 5'h6 : _GEN_7046; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7060 = 2'h1 == opidx ? 5'h6 : _GEN_7047; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7061 = 2'h2 == opidx ? 5'h6 : _GEN_7048; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7062 = 2'h3 == opidx ? 5'h6 : _GEN_7049; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7063 = 2'h0 == opidx ? regback_1 : _GEN_7050; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7064 = 2'h1 == opidx ? regback_1 : _GEN_7051; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7065 = 2'h2 == opidx ? regback_1 : _GEN_7052; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7066 = 2'h3 == opidx ? regback_1 : _GEN_7053; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7067 = ~_GEN_1128 ? _cnt_T : _GEN_7054; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7068 = cnt[33] ? _GEN_7055 : _GEN_7042; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7069 = cnt[33] ? _GEN_7056 : _GEN_7043; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7070 = cnt[33] ? _GEN_7057 : _GEN_7044; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7071 = cnt[33] ? _GEN_7058 : _GEN_7045; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7072 = cnt[33] ? _GEN_7059 : _GEN_7046; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7073 = cnt[33] ? _GEN_7060 : _GEN_7047; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7074 = cnt[33] ? _GEN_7061 : _GEN_7048; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7075 = cnt[33] ? _GEN_7062 : _GEN_7049; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7076 = cnt[33] ? _GEN_7063 : _GEN_7050; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7077 = cnt[33] ? _GEN_7064 : _GEN_7051; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7078 = cnt[33] ? _GEN_7065 : _GEN_7052; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7079 = cnt[33] ? _GEN_7066 : _GEN_7053; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7080 = cnt[33] ? _GEN_7067 : _GEN_7054; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7081 = _GEN_145 | _GEN_7068; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7082 = _GEN_146 | _GEN_7069; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7083 = _GEN_147 | _GEN_7070; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7084 = _GEN_148 | _GEN_7071; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7085 = 2'h0 == opidx ? 5'h7 : _GEN_7072; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7086 = 2'h1 == opidx ? 5'h7 : _GEN_7073; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7087 = 2'h2 == opidx ? 5'h7 : _GEN_7074; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7088 = 2'h3 == opidx ? 5'h7 : _GEN_7075; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7089 = 2'h0 == opidx ? regback_2 : _GEN_7076; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7090 = 2'h1 == opidx ? regback_2 : _GEN_7077; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7091 = 2'h2 == opidx ? regback_2 : _GEN_7078; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7092 = 2'h3 == opidx ? regback_2 : _GEN_7079; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7093 = ~_GEN_1128 ? _cnt_T : _GEN_7080; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7094 = cnt[34] ? _GEN_7081 : _GEN_7068; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7095 = cnt[34] ? _GEN_7082 : _GEN_7069; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7096 = cnt[34] ? _GEN_7083 : _GEN_7070; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7097 = cnt[34] ? _GEN_7084 : _GEN_7071; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7098 = cnt[34] ? _GEN_7085 : _GEN_7072; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7099 = cnt[34] ? _GEN_7086 : _GEN_7073; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7100 = cnt[34] ? _GEN_7087 : _GEN_7074; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7101 = cnt[34] ? _GEN_7088 : _GEN_7075; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7102 = cnt[34] ? _GEN_7089 : _GEN_7076; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7103 = cnt[34] ? _GEN_7090 : _GEN_7077; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7104 = cnt[34] ? _GEN_7091 : _GEN_7078; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7105 = cnt[34] ? _GEN_7092 : _GEN_7079; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7106 = cnt[34] ? _GEN_7093 : _GEN_7080; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7107 = _GEN_145 | _GEN_7094; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7108 = _GEN_146 | _GEN_7095; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7109 = _GEN_147 | _GEN_7096; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7110 = _GEN_148 | _GEN_7097; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7111 = 2'h0 == opidx ? 5'h8 : _GEN_7098; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7112 = 2'h1 == opidx ? 5'h8 : _GEN_7099; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7113 = 2'h2 == opidx ? 5'h8 : _GEN_7100; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7114 = 2'h3 == opidx ? 5'h8 : _GEN_7101; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7115 = 2'h0 == opidx ? regback_3 : _GEN_7102; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7116 = 2'h1 == opidx ? regback_3 : _GEN_7103; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7117 = 2'h2 == opidx ? regback_3 : _GEN_7104; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7118 = 2'h3 == opidx ? regback_3 : _GEN_7105; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7119 = ~_GEN_1128 ? _cnt_T : _GEN_7106; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7120 = cnt[35] ? _GEN_7107 : _GEN_7094; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7121 = cnt[35] ? _GEN_7108 : _GEN_7095; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7122 = cnt[35] ? _GEN_7109 : _GEN_7096; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7123 = cnt[35] ? _GEN_7110 : _GEN_7097; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7124 = cnt[35] ? _GEN_7111 : _GEN_7098; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7125 = cnt[35] ? _GEN_7112 : _GEN_7099; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7126 = cnt[35] ? _GEN_7113 : _GEN_7100; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7127 = cnt[35] ? _GEN_7114 : _GEN_7101; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7128 = cnt[35] ? _GEN_7115 : _GEN_7102; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7129 = cnt[35] ? _GEN_7116 : _GEN_7103; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7130 = cnt[35] ? _GEN_7117 : _GEN_7104; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7131 = cnt[35] ? _GEN_7118 : _GEN_7105; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7132 = cnt[35] ? _GEN_7119 : _GEN_7106; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7133 = _GEN_145 | _GEN_7120; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7134 = _GEN_146 | _GEN_7121; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7135 = _GEN_147 | _GEN_7122; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7136 = _GEN_148 | _GEN_7123; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7137 = 2'h0 == opidx ? 5'h9 : _GEN_7124; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7138 = 2'h1 == opidx ? 5'h9 : _GEN_7125; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7139 = 2'h2 == opidx ? 5'h9 : _GEN_7126; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7140 = 2'h3 == opidx ? 5'h9 : _GEN_7127; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7141 = 2'h0 == opidx ? regback_4 : _GEN_7128; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7142 = 2'h1 == opidx ? regback_4 : _GEN_7129; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7143 = 2'h2 == opidx ? regback_4 : _GEN_7130; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7144 = 2'h3 == opidx ? regback_4 : _GEN_7131; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7145 = ~_GEN_1128 ? _cnt_T : _GEN_7132; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7146 = cnt[36] ? _GEN_7133 : _GEN_7120; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7147 = cnt[36] ? _GEN_7134 : _GEN_7121; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7148 = cnt[36] ? _GEN_7135 : _GEN_7122; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7149 = cnt[36] ? _GEN_7136 : _GEN_7123; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7150 = cnt[36] ? _GEN_7137 : _GEN_7124; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7151 = cnt[36] ? _GEN_7138 : _GEN_7125; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7152 = cnt[36] ? _GEN_7139 : _GEN_7126; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7153 = cnt[36] ? _GEN_7140 : _GEN_7127; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7154 = cnt[36] ? _GEN_7141 : _GEN_7128; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7155 = cnt[36] ? _GEN_7142 : _GEN_7129; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7156 = cnt[36] ? _GEN_7143 : _GEN_7130; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7157 = cnt[36] ? _GEN_7144 : _GEN_7131; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7158 = cnt[36] ? _GEN_7145 : _GEN_7132; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7159 = _GEN_145 | _GEN_7146; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7160 = _GEN_146 | _GEN_7147; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7161 = _GEN_147 | _GEN_7148; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7162 = _GEN_148 | _GEN_7149; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7163 = 2'h0 == opidx ? 5'ha : _GEN_7150; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7164 = 2'h1 == opidx ? 5'ha : _GEN_7151; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7165 = 2'h2 == opidx ? 5'ha : _GEN_7152; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7166 = 2'h3 == opidx ? 5'ha : _GEN_7153; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7167 = 2'h0 == opidx ? regback_5 : _GEN_7154; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7168 = 2'h1 == opidx ? regback_5 : _GEN_7155; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7169 = 2'h2 == opidx ? regback_5 : _GEN_7156; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7170 = 2'h3 == opidx ? regback_5 : _GEN_7157; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7171 = ~_GEN_1128 ? _cnt_T : _GEN_7158; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7172 = cnt[37] ? _GEN_7159 : _GEN_7146; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7173 = cnt[37] ? _GEN_7160 : _GEN_7147; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7174 = cnt[37] ? _GEN_7161 : _GEN_7148; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7175 = cnt[37] ? _GEN_7162 : _GEN_7149; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7176 = cnt[37] ? _GEN_7163 : _GEN_7150; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7177 = cnt[37] ? _GEN_7164 : _GEN_7151; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7178 = cnt[37] ? _GEN_7165 : _GEN_7152; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7179 = cnt[37] ? _GEN_7166 : _GEN_7153; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7180 = cnt[37] ? _GEN_7167 : _GEN_7154; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7181 = cnt[37] ? _GEN_7168 : _GEN_7155; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7182 = cnt[37] ? _GEN_7169 : _GEN_7156; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7183 = cnt[37] ? _GEN_7170 : _GEN_7157; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7184 = cnt[37] ? _GEN_7171 : _GEN_7158; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7185 = _GEN_145 | _GEN_7172; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7186 = _GEN_146 | _GEN_7173; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7187 = _GEN_147 | _GEN_7174; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7188 = _GEN_148 | _GEN_7175; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7189 = 2'h0 == opidx ? 5'hb : _GEN_7176; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7190 = 2'h1 == opidx ? 5'hb : _GEN_7177; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7191 = 2'h2 == opidx ? 5'hb : _GEN_7178; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7192 = 2'h3 == opidx ? 5'hb : _GEN_7179; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7193 = 2'h0 == opidx ? regback_6 : _GEN_7180; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7194 = 2'h1 == opidx ? regback_6 : _GEN_7181; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7195 = 2'h2 == opidx ? regback_6 : _GEN_7182; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7196 = 2'h3 == opidx ? regback_6 : _GEN_7183; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7197 = ~_GEN_1128 ? _cnt_T : _GEN_7184; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7198 = cnt[38] ? _GEN_7185 : _GEN_7172; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7199 = cnt[38] ? _GEN_7186 : _GEN_7173; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7200 = cnt[38] ? _GEN_7187 : _GEN_7174; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7201 = cnt[38] ? _GEN_7188 : _GEN_7175; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7202 = cnt[38] ? _GEN_7189 : _GEN_7176; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7203 = cnt[38] ? _GEN_7190 : _GEN_7177; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7204 = cnt[38] ? _GEN_7191 : _GEN_7178; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7205 = cnt[38] ? _GEN_7192 : _GEN_7179; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7206 = cnt[38] ? _GEN_7193 : _GEN_7180; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7207 = cnt[38] ? _GEN_7194 : _GEN_7181; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7208 = cnt[38] ? _GEN_7195 : _GEN_7182; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7209 = cnt[38] ? _GEN_7196 : _GEN_7183; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7210 = cnt[38] ? _GEN_7197 : _GEN_7184; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7211 = _GEN_145 | _GEN_7198; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7212 = _GEN_146 | _GEN_7199; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7213 = _GEN_147 | _GEN_7200; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7214 = _GEN_148 | _GEN_7201; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7215 = 2'h0 == opidx ? 5'hc : _GEN_7202; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7216 = 2'h1 == opidx ? 5'hc : _GEN_7203; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7217 = 2'h2 == opidx ? 5'hc : _GEN_7204; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7218 = 2'h3 == opidx ? 5'hc : _GEN_7205; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7219 = 2'h0 == opidx ? regback_7 : _GEN_7206; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7220 = 2'h1 == opidx ? regback_7 : _GEN_7207; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7221 = 2'h2 == opidx ? regback_7 : _GEN_7208; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7222 = 2'h3 == opidx ? regback_7 : _GEN_7209; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7223 = ~_GEN_1128 ? _cnt_T : _GEN_7210; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7224 = cnt[39] ? _GEN_7211 : _GEN_7198; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7225 = cnt[39] ? _GEN_7212 : _GEN_7199; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7226 = cnt[39] ? _GEN_7213 : _GEN_7200; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7227 = cnt[39] ? _GEN_7214 : _GEN_7201; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7228 = cnt[39] ? _GEN_7215 : _GEN_7202; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7229 = cnt[39] ? _GEN_7216 : _GEN_7203; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7230 = cnt[39] ? _GEN_7217 : _GEN_7204; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7231 = cnt[39] ? _GEN_7218 : _GEN_7205; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7232 = cnt[39] ? _GEN_7219 : _GEN_7206; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7233 = cnt[39] ? _GEN_7220 : _GEN_7207; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7234 = cnt[39] ? _GEN_7221 : _GEN_7208; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7235 = cnt[39] ? _GEN_7222 : _GEN_7209; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7236 = cnt[39] ? _GEN_7223 : _GEN_7210; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7237 = _GEN_145 | _GEN_7224; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7238 = _GEN_146 | _GEN_7225; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7239 = _GEN_147 | _GEN_7226; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7240 = _GEN_148 | _GEN_7227; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7241 = 2'h0 == opidx ? 5'hd : _GEN_7228; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7242 = 2'h1 == opidx ? 5'hd : _GEN_7229; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7243 = 2'h2 == opidx ? 5'hd : _GEN_7230; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7244 = 2'h3 == opidx ? 5'hd : _GEN_7231; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7245 = 2'h0 == opidx ? regback_8 : _GEN_7232; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7246 = 2'h1 == opidx ? regback_8 : _GEN_7233; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7247 = 2'h2 == opidx ? regback_8 : _GEN_7234; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7248 = 2'h3 == opidx ? regback_8 : _GEN_7235; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7249 = ~_GEN_1128 ? _cnt_T : _GEN_7236; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7250 = cnt[40] ? _GEN_7237 : _GEN_7224; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7251 = cnt[40] ? _GEN_7238 : _GEN_7225; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7252 = cnt[40] ? _GEN_7239 : _GEN_7226; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_7253 = cnt[40] ? _GEN_7240 : _GEN_7227; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7254 = cnt[40] ? _GEN_7241 : _GEN_7228; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7255 = cnt[40] ? _GEN_7242 : _GEN_7229; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7256 = cnt[40] ? _GEN_7243 : _GEN_7230; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_7257 = cnt[40] ? _GEN_7244 : _GEN_7231; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7258 = cnt[40] ? _GEN_7245 : _GEN_7232; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7259 = cnt[40] ? _GEN_7246 : _GEN_7233; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7260 = cnt[40] ? _GEN_7247 : _GEN_7234; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_7261 = cnt[40] ? _GEN_7248 : _GEN_7235; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7262 = cnt[40] ? _GEN_7249 : _GEN_7236; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_7263 = pgbuf_cpu_pos == pgbuf_uart_pos ? 129'h1 : _GEN_7262; // @[NulCtrlMP.scala 857:52 858:21]
  wire [4:0] _GEN_7264 = pgbuf_cpu_pos == pgbuf_uart_pos ? 5'h1f : _GEN_4935; // @[NulCtrlMP.scala 857:52 859:23]
  wire [11:0] _GEN_7265 = pgbuf_cpu_pos == pgbuf_uart_pos ? 12'h0 : _GEN_7000; // @[NulCtrlMP.scala 857:52 860:31]
  wire [11:0] _GEN_7266 = pgbuf_cpu_pos == pgbuf_uart_pos ? 12'h0 : pgbuf_uart_pos; // @[NulCtrlMP.scala 857:52 861:32 819:33]
  wire [128:0] _GEN_7267 = cnt[41] ? _GEN_7263 : _GEN_7262; // @[NulCtrlMP.scala 856:23]
  wire [4:0] _GEN_7268 = cnt[41] ? _GEN_7264 : _GEN_4935; // @[NulCtrlMP.scala 856:23]
  wire [11:0] _GEN_7269 = cnt[41] ? _GEN_7265 : _GEN_7000; // @[NulCtrlMP.scala 856:23]
  wire [11:0] _GEN_7270 = cnt[41] ? _GEN_7266 : pgbuf_uart_pos; // @[NulCtrlMP.scala 856:23 819:33]
  wire [6:0] shift = pgbuf_uart_pos[2:0] * 4'h8; // @[NulCtrlMP.scala 868:46]
  wire [63:0] _GEN_7272 = 6'h1 == pgbuf_uart_pos[8:3] ? pgbuf_div8_1 : pgbuf_div8_0; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7273 = 6'h2 == pgbuf_uart_pos[8:3] ? pgbuf_div8_2 : _GEN_7272; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7274 = 6'h3 == pgbuf_uart_pos[8:3] ? pgbuf_div8_3 : _GEN_7273; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7275 = 6'h4 == pgbuf_uart_pos[8:3] ? pgbuf_div8_4 : _GEN_7274; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7276 = 6'h5 == pgbuf_uart_pos[8:3] ? pgbuf_div8_5 : _GEN_7275; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7277 = 6'h6 == pgbuf_uart_pos[8:3] ? pgbuf_div8_6 : _GEN_7276; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7278 = 6'h7 == pgbuf_uart_pos[8:3] ? pgbuf_div8_7 : _GEN_7277; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7279 = 6'h8 == pgbuf_uart_pos[8:3] ? pgbuf_div8_8 : _GEN_7278; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7280 = 6'h9 == pgbuf_uart_pos[8:3] ? pgbuf_div8_9 : _GEN_7279; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7281 = 6'ha == pgbuf_uart_pos[8:3] ? pgbuf_div8_10 : _GEN_7280; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7282 = 6'hb == pgbuf_uart_pos[8:3] ? pgbuf_div8_11 : _GEN_7281; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7283 = 6'hc == pgbuf_uart_pos[8:3] ? pgbuf_div8_12 : _GEN_7282; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7284 = 6'hd == pgbuf_uart_pos[8:3] ? pgbuf_div8_13 : _GEN_7283; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7285 = 6'he == pgbuf_uart_pos[8:3] ? pgbuf_div8_14 : _GEN_7284; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7286 = 6'hf == pgbuf_uart_pos[8:3] ? pgbuf_div8_15 : _GEN_7285; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7287 = 6'h10 == pgbuf_uart_pos[8:3] ? pgbuf_div8_16 : _GEN_7286; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7288 = 6'h11 == pgbuf_uart_pos[8:3] ? pgbuf_div8_17 : _GEN_7287; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7289 = 6'h12 == pgbuf_uart_pos[8:3] ? pgbuf_div8_18 : _GEN_7288; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7290 = 6'h13 == pgbuf_uart_pos[8:3] ? pgbuf_div8_19 : _GEN_7289; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7291 = 6'h14 == pgbuf_uart_pos[8:3] ? pgbuf_div8_20 : _GEN_7290; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7292 = 6'h15 == pgbuf_uart_pos[8:3] ? pgbuf_div8_21 : _GEN_7291; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7293 = 6'h16 == pgbuf_uart_pos[8:3] ? pgbuf_div8_22 : _GEN_7292; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7294 = 6'h17 == pgbuf_uart_pos[8:3] ? pgbuf_div8_23 : _GEN_7293; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7295 = 6'h18 == pgbuf_uart_pos[8:3] ? pgbuf_div8_24 : _GEN_7294; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7296 = 6'h19 == pgbuf_uart_pos[8:3] ? pgbuf_div8_25 : _GEN_7295; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7297 = 6'h1a == pgbuf_uart_pos[8:3] ? pgbuf_div8_26 : _GEN_7296; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7298 = 6'h1b == pgbuf_uart_pos[8:3] ? pgbuf_div8_27 : _GEN_7297; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7299 = 6'h1c == pgbuf_uart_pos[8:3] ? pgbuf_div8_28 : _GEN_7298; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7300 = 6'h1d == pgbuf_uart_pos[8:3] ? pgbuf_div8_29 : _GEN_7299; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7301 = 6'h1e == pgbuf_uart_pos[8:3] ? pgbuf_div8_30 : _GEN_7300; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7302 = 6'h1f == pgbuf_uart_pos[8:3] ? pgbuf_div8_31 : _GEN_7301; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7303 = 6'h20 == pgbuf_uart_pos[8:3] ? pgbuf_div8_32 : _GEN_7302; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7304 = 6'h21 == pgbuf_uart_pos[8:3] ? pgbuf_div8_33 : _GEN_7303; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7305 = 6'h22 == pgbuf_uart_pos[8:3] ? pgbuf_div8_34 : _GEN_7304; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7306 = 6'h23 == pgbuf_uart_pos[8:3] ? pgbuf_div8_35 : _GEN_7305; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7307 = 6'h24 == pgbuf_uart_pos[8:3] ? pgbuf_div8_36 : _GEN_7306; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7308 = 6'h25 == pgbuf_uart_pos[8:3] ? pgbuf_div8_37 : _GEN_7307; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7309 = 6'h26 == pgbuf_uart_pos[8:3] ? pgbuf_div8_38 : _GEN_7308; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7310 = 6'h27 == pgbuf_uart_pos[8:3] ? pgbuf_div8_39 : _GEN_7309; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7311 = 6'h28 == pgbuf_uart_pos[8:3] ? pgbuf_div8_40 : _GEN_7310; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7312 = 6'h29 == pgbuf_uart_pos[8:3] ? pgbuf_div8_41 : _GEN_7311; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7313 = 6'h2a == pgbuf_uart_pos[8:3] ? pgbuf_div8_42 : _GEN_7312; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7314 = 6'h2b == pgbuf_uart_pos[8:3] ? pgbuf_div8_43 : _GEN_7313; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7315 = 6'h2c == pgbuf_uart_pos[8:3] ? pgbuf_div8_44 : _GEN_7314; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7316 = 6'h2d == pgbuf_uart_pos[8:3] ? pgbuf_div8_45 : _GEN_7315; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7317 = 6'h2e == pgbuf_uart_pos[8:3] ? pgbuf_div8_46 : _GEN_7316; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7318 = 6'h2f == pgbuf_uart_pos[8:3] ? pgbuf_div8_47 : _GEN_7317; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7319 = 6'h30 == pgbuf_uart_pos[8:3] ? pgbuf_div8_48 : _GEN_7318; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7320 = 6'h31 == pgbuf_uart_pos[8:3] ? pgbuf_div8_49 : _GEN_7319; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7321 = 6'h32 == pgbuf_uart_pos[8:3] ? pgbuf_div8_50 : _GEN_7320; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7322 = 6'h33 == pgbuf_uart_pos[8:3] ? pgbuf_div8_51 : _GEN_7321; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7323 = 6'h34 == pgbuf_uart_pos[8:3] ? pgbuf_div8_52 : _GEN_7322; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7324 = 6'h35 == pgbuf_uart_pos[8:3] ? pgbuf_div8_53 : _GEN_7323; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7325 = 6'h36 == pgbuf_uart_pos[8:3] ? pgbuf_div8_54 : _GEN_7324; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7326 = 6'h37 == pgbuf_uart_pos[8:3] ? pgbuf_div8_55 : _GEN_7325; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7327 = 6'h38 == pgbuf_uart_pos[8:3] ? pgbuf_div8_56 : _GEN_7326; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7328 = 6'h39 == pgbuf_uart_pos[8:3] ? pgbuf_div8_57 : _GEN_7327; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7329 = 6'h3a == pgbuf_uart_pos[8:3] ? pgbuf_div8_58 : _GEN_7328; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7330 = 6'h3b == pgbuf_uart_pos[8:3] ? pgbuf_div8_59 : _GEN_7329; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7331 = 6'h3c == pgbuf_uart_pos[8:3] ? pgbuf_div8_60 : _GEN_7330; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7332 = 6'h3d == pgbuf_uart_pos[8:3] ? pgbuf_div8_61 : _GEN_7331; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7333 = 6'h3e == pgbuf_uart_pos[8:3] ? pgbuf_div8_62 : _GEN_7332; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _GEN_7334 = 6'h3f == pgbuf_uart_pos[8:3] ? pgbuf_div8_63 : _GEN_7333; // @[NulCtrlMP.scala 869:{33,33}]
  wire [63:0] _io_tx_bits_T_3 = _GEN_7334 >> shift; // @[NulCtrlMP.scala 869:33]
  wire [11:0] _pgbuf_uart_pos_T_1 = pgbuf_uart_pos + 12'h1; // @[NulCtrlMP.scala 871:50]
  wire [11:0] _GEN_7335 = io_tx_ready ? _pgbuf_uart_pos_T_1 : _GEN_7270; // @[NulCtrlMP.scala 870:31 871:32]
  wire  _GEN_7336 = cnt[9:0] == 10'h0 & pgbuf_cpu_pos > pgbuf_uart_pos | _GEN_5117; // @[NulCtrlMP.scala 865:67 866:25]
  wire [7:0] _GEN_7337 = cnt[9:0] == 10'h0 & pgbuf_cpu_pos > pgbuf_uart_pos ? _io_tx_bits_T_3[7:0] : _GEN_5118; // @[NulCtrlMP.scala 865:67 869:24]
  wire [11:0] _GEN_7338 = cnt[9:0] == 10'h0 & pgbuf_cpu_pos > pgbuf_uart_pos ? _GEN_7335 : _GEN_7270; // @[NulCtrlMP.scala 865:67]
  wire  _GEN_7339 = state == 5'h12 ? _GEN_6925 : _GEN_4895; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7340 = state == 5'h12 ? _GEN_6926 : _GEN_4896; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7341 = state == 5'h12 ? _GEN_6927 : _GEN_4897; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7342 = state == 5'h12 ? _GEN_6928 : _GEN_4898; // @[NulCtrlMP.scala 822:32]
  wire [4:0] _GEN_7343 = state == 5'h12 ? _GEN_7254 : _GEN_4899; // @[NulCtrlMP.scala 822:32]
  wire [4:0] _GEN_7344 = state == 5'h12 ? _GEN_7255 : _GEN_4900; // @[NulCtrlMP.scala 822:32]
  wire [4:0] _GEN_7345 = state == 5'h12 ? _GEN_7256 : _GEN_4901; // @[NulCtrlMP.scala 822:32]
  wire [4:0] _GEN_7346 = state == 5'h12 ? _GEN_7257 : _GEN_4902; // @[NulCtrlMP.scala 822:32]
  wire [128:0] _GEN_7347 = state == 5'h12 ? _GEN_7267 : _GEN_4903; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7348 = state == 5'h12 ? _GEN_4955 : _GEN_4904; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7349 = state == 5'h12 ? _GEN_4975 : _GEN_4905; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7350 = state == 5'h12 ? _GEN_4995 : _GEN_4906; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7351 = state == 5'h12 ? _GEN_5015 : _GEN_4907; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7352 = state == 5'h12 ? _GEN_5035 : _GEN_4908; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7353 = state == 5'h12 ? _GEN_5055 : _GEN_4909; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7354 = state == 5'h12 ? _GEN_5075 : _GEN_4910; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7355 = state == 5'h12 ? _GEN_5095 : _GEN_4911; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7356 = state == 5'h12 ? _GEN_5115 : _GEN_4912; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7357 = state == 5'h12 ? _GEN_7336 : _GEN_1102; // @[NulCtrlMP.scala 822:32]
  wire [7:0] _GEN_7358 = state == 5'h12 ? _GEN_7337 : _GEN_1103; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7359 = state == 5'h12 ? _GEN_7250 : _GEN_4914; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7360 = state == 5'h12 ? _GEN_7251 : _GEN_4915; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7361 = state == 5'h12 ? _GEN_7252 : _GEN_4916; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7362 = state == 5'h12 ? _GEN_7253 : _GEN_4917; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7363 = state == 5'h12 ? _GEN_7258 : _GEN_4918; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7364 = state == 5'h12 ? _GEN_7259 : _GEN_4919; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7365 = state == 5'h12 ? _GEN_7260 : _GEN_4920; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7366 = state == 5'h12 ? _GEN_7261 : _GEN_4921; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7367 = state == 5'h12 ? _GEN_7010 : _GEN_4922; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7368 = state == 5'h12 ? _GEN_7011 : _GEN_4923; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7369 = state == 5'h12 ? _GEN_7012 : _GEN_4924; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7370 = state == 5'h12 ? _GEN_7013 : _GEN_4925; // @[NulCtrlMP.scala 822:32]
  wire [31:0] _GEN_7371 = state == 5'h12 ? _GEN_7014 : _GEN_4926; // @[NulCtrlMP.scala 822:32]
  wire [31:0] _GEN_7372 = state == 5'h12 ? _GEN_7015 : _GEN_4927; // @[NulCtrlMP.scala 822:32]
  wire [31:0] _GEN_7373 = state == 5'h12 ? _GEN_7016 : _GEN_4928; // @[NulCtrlMP.scala 822:32]
  wire [31:0] _GEN_7374 = state == 5'h12 ? _GEN_7017 : _GEN_4929; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7375 = state == 5'h12 ? _GEN_7024 : _GEN_4930; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7376 = state == 5'h12 ? _GEN_7025 : _GEN_4931; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7377 = state == 5'h12 ? _GEN_7026 : _GEN_4932; // @[NulCtrlMP.scala 822:32]
  wire  _GEN_7378 = state == 5'h12 ? _GEN_7027 : _GEN_4933; // @[NulCtrlMP.scala 822:32]
  wire [63:0] _GEN_7379 = state == 5'h12 ? _GEN_6934 : pgbuf_div8_0; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7380 = state == 5'h12 ? _GEN_6935 : pgbuf_div8_1; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7381 = state == 5'h12 ? _GEN_6936 : pgbuf_div8_2; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7382 = state == 5'h12 ? _GEN_6937 : pgbuf_div8_3; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7383 = state == 5'h12 ? _GEN_6938 : pgbuf_div8_4; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7384 = state == 5'h12 ? _GEN_6939 : pgbuf_div8_5; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7385 = state == 5'h12 ? _GEN_6940 : pgbuf_div8_6; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7386 = state == 5'h12 ? _GEN_6941 : pgbuf_div8_7; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7387 = state == 5'h12 ? _GEN_6942 : pgbuf_div8_8; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7388 = state == 5'h12 ? _GEN_6943 : pgbuf_div8_9; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7389 = state == 5'h12 ? _GEN_6944 : pgbuf_div8_10; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7390 = state == 5'h12 ? _GEN_6945 : pgbuf_div8_11; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7391 = state == 5'h12 ? _GEN_6946 : pgbuf_div8_12; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7392 = state == 5'h12 ? _GEN_6947 : pgbuf_div8_13; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7393 = state == 5'h12 ? _GEN_6948 : pgbuf_div8_14; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7394 = state == 5'h12 ? _GEN_6949 : pgbuf_div8_15; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7395 = state == 5'h12 ? _GEN_6950 : pgbuf_div8_16; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7396 = state == 5'h12 ? _GEN_6951 : pgbuf_div8_17; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7397 = state == 5'h12 ? _GEN_6952 : pgbuf_div8_18; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7398 = state == 5'h12 ? _GEN_6953 : pgbuf_div8_19; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7399 = state == 5'h12 ? _GEN_6954 : pgbuf_div8_20; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7400 = state == 5'h12 ? _GEN_6955 : pgbuf_div8_21; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7401 = state == 5'h12 ? _GEN_6956 : pgbuf_div8_22; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7402 = state == 5'h12 ? _GEN_6957 : pgbuf_div8_23; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7403 = state == 5'h12 ? _GEN_6958 : pgbuf_div8_24; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7404 = state == 5'h12 ? _GEN_6959 : pgbuf_div8_25; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7405 = state == 5'h12 ? _GEN_6960 : pgbuf_div8_26; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7406 = state == 5'h12 ? _GEN_6961 : pgbuf_div8_27; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7407 = state == 5'h12 ? _GEN_6962 : pgbuf_div8_28; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7408 = state == 5'h12 ? _GEN_6963 : pgbuf_div8_29; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7409 = state == 5'h12 ? _GEN_6964 : pgbuf_div8_30; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7410 = state == 5'h12 ? _GEN_6965 : pgbuf_div8_31; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7411 = state == 5'h12 ? _GEN_6966 : pgbuf_div8_32; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7412 = state == 5'h12 ? _GEN_6967 : pgbuf_div8_33; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7413 = state == 5'h12 ? _GEN_6968 : pgbuf_div8_34; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7414 = state == 5'h12 ? _GEN_6969 : pgbuf_div8_35; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7415 = state == 5'h12 ? _GEN_6970 : pgbuf_div8_36; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7416 = state == 5'h12 ? _GEN_6971 : pgbuf_div8_37; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7417 = state == 5'h12 ? _GEN_6972 : pgbuf_div8_38; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7418 = state == 5'h12 ? _GEN_6973 : pgbuf_div8_39; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7419 = state == 5'h12 ? _GEN_6974 : pgbuf_div8_40; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7420 = state == 5'h12 ? _GEN_6975 : pgbuf_div8_41; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7421 = state == 5'h12 ? _GEN_6976 : pgbuf_div8_42; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7422 = state == 5'h12 ? _GEN_6977 : pgbuf_div8_43; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7423 = state == 5'h12 ? _GEN_6978 : pgbuf_div8_44; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7424 = state == 5'h12 ? _GEN_6979 : pgbuf_div8_45; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7425 = state == 5'h12 ? _GEN_6980 : pgbuf_div8_46; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7426 = state == 5'h12 ? _GEN_6981 : pgbuf_div8_47; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7427 = state == 5'h12 ? _GEN_6982 : pgbuf_div8_48; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7428 = state == 5'h12 ? _GEN_6983 : pgbuf_div8_49; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7429 = state == 5'h12 ? _GEN_6984 : pgbuf_div8_50; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7430 = state == 5'h12 ? _GEN_6985 : pgbuf_div8_51; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7431 = state == 5'h12 ? _GEN_6986 : pgbuf_div8_52; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7432 = state == 5'h12 ? _GEN_6987 : pgbuf_div8_53; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7433 = state == 5'h12 ? _GEN_6988 : pgbuf_div8_54; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7434 = state == 5'h12 ? _GEN_6989 : pgbuf_div8_55; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7435 = state == 5'h12 ? _GEN_6990 : pgbuf_div8_56; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7436 = state == 5'h12 ? _GEN_6991 : pgbuf_div8_57; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7437 = state == 5'h12 ? _GEN_6992 : pgbuf_div8_58; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7438 = state == 5'h12 ? _GEN_6993 : pgbuf_div8_59; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7439 = state == 5'h12 ? _GEN_6994 : pgbuf_div8_60; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7440 = state == 5'h12 ? _GEN_6995 : pgbuf_div8_61; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7441 = state == 5'h12 ? _GEN_6996 : pgbuf_div8_62; // @[NulCtrlMP.scala 818:29 822:32]
  wire [63:0] _GEN_7442 = state == 5'h12 ? _GEN_6997 : pgbuf_div8_63; // @[NulCtrlMP.scala 818:29 822:32]
  wire [11:0] _GEN_7443 = state == 5'h12 ? _GEN_7269 : pgbuf_cpu_pos; // @[NulCtrlMP.scala 820:32 822:32]
  wire [4:0] _GEN_7444 = state == 5'h12 ? _GEN_7268 : _GEN_4935; // @[NulCtrlMP.scala 822:32]
  wire [11:0] _GEN_7445 = state == 5'h12 ? _GEN_7338 : pgbuf_uart_pos; // @[NulCtrlMP.scala 822:32 819:33]
  reg [3:0] wt_byte_cnt; // @[NulCtrlMP.scala 876:30]
  reg [7:0] wt_byte_buf_0; // @[NulCtrlMP.scala 877:30]
  reg [7:0] wt_byte_buf_1; // @[NulCtrlMP.scala 877:30]
  reg [7:0] wt_byte_buf_2; // @[NulCtrlMP.scala 877:30]
  reg [7:0] wt_byte_buf_3; // @[NulCtrlMP.scala 877:30]
  reg [7:0] wt_byte_buf_4; // @[NulCtrlMP.scala 877:30]
  reg [7:0] wt_byte_buf_5; // @[NulCtrlMP.scala 877:30]
  reg [7:0] wt_byte_buf_6; // @[NulCtrlMP.scala 877:30]
  wire  _T_555 = pgbuf_uart_pos != 12'h200; // @[NulCtrlMP.scala 880:29]
  wire  _GEN_7446 = pgbuf_uart_pos != 12'h200 | _GEN_125; // @[NulCtrlMP.scala 880:40 881:25]
  wire [63:0] _pgbuf_div8_T = {io_rx_bits,wt_byte_buf_6,wt_byte_buf_5,wt_byte_buf_4,wt_byte_buf_3,wt_byte_buf_2,
    wt_byte_buf_1,wt_byte_buf_0}; // @[Cat.scala 31:58]
  wire [63:0] _GEN_7455 = 6'h0 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7379; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7456 = 6'h1 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7380; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7457 = 6'h2 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7381; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7458 = 6'h3 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7382; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7459 = 6'h4 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7383; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7460 = 6'h5 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7384; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7461 = 6'h6 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7385; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7462 = 6'h7 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7386; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7463 = 6'h8 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7387; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7464 = 6'h9 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7388; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7465 = 6'ha == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7389; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7466 = 6'hb == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7390; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7467 = 6'hc == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7391; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7468 = 6'hd == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7392; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7469 = 6'he == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7393; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7470 = 6'hf == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7394; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7471 = 6'h10 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7395; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7472 = 6'h11 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7396; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7473 = 6'h12 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7397; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7474 = 6'h13 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7398; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7475 = 6'h14 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7399; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7476 = 6'h15 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7400; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7477 = 6'h16 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7401; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7478 = 6'h17 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7402; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7479 = 6'h18 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7403; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7480 = 6'h19 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7404; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7481 = 6'h1a == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7405; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7482 = 6'h1b == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7406; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7483 = 6'h1c == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7407; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7484 = 6'h1d == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7408; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7485 = 6'h1e == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7409; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7486 = 6'h1f == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7410; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7487 = 6'h20 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7411; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7488 = 6'h21 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7412; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7489 = 6'h22 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7413; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7490 = 6'h23 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7414; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7491 = 6'h24 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7415; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7492 = 6'h25 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7416; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7493 = 6'h26 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7417; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7494 = 6'h27 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7418; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7495 = 6'h28 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7419; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7496 = 6'h29 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7420; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7497 = 6'h2a == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7421; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7498 = 6'h2b == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7422; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7499 = 6'h2c == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7423; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7500 = 6'h2d == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7424; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7501 = 6'h2e == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7425; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7502 = 6'h2f == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7426; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7503 = 6'h30 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7427; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7504 = 6'h31 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7428; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7505 = 6'h32 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7429; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7506 = 6'h33 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7430; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7507 = 6'h34 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7431; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7508 = 6'h35 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7432; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7509 = 6'h36 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7433; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7510 = 6'h37 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7434; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7511 = 6'h38 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7435; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7512 = 6'h39 == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7436; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7513 = 6'h3a == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7437; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7514 = 6'h3b == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7438; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7515 = 6'h3c == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7439; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7516 = 6'h3d == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7440; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7517 = 6'h3e == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7441; // @[NulCtrlMP.scala 887:{49,49}]
  wire [63:0] _GEN_7518 = 6'h3f == pgbuf_uart_pos[8:3] ? _pgbuf_div8_T : _GEN_7442; // @[NulCtrlMP.scala 887:{49,49}]
  wire [11:0] _pgbuf_uart_pos_T_3 = pgbuf_uart_pos + 12'h8; // @[NulCtrlMP.scala 888:50]
  wire [3:0] _wt_byte_cnt_T_1 = wt_byte_cnt + 4'h1; // @[NulCtrlMP.scala 890:44]
  wire [3:0] _GEN_7519 = wt_byte_cnt == 4'h7 ? 4'h0 : _wt_byte_cnt_T_1; // @[NulCtrlMP.scala 885:39 886:29 890:29]
  wire [11:0] _GEN_7584 = wt_byte_cnt == 4'h7 ? _pgbuf_uart_pos_T_3 : _GEN_7445; // @[NulCtrlMP.scala 885:39 888:32]
  wire  _GEN_7659 = _GEN_145 | _GEN_7339; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7660 = _GEN_146 | _GEN_7340; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7661 = _GEN_147 | _GEN_7341; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7662 = _GEN_148 | _GEN_7342; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_7663 = 2'h0 == opidx ? 5'h5 : _GEN_7343; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7664 = 2'h1 == opidx ? 5'h5 : _GEN_7344; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7665 = 2'h2 == opidx ? 5'h5 : _GEN_7345; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7666 = 2'h3 == opidx ? 5'h5 : _GEN_7346; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_7667 = _T_122 ? _cnt_T : _GEN_7347; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_7669 = cnt[0] ? _GEN_7659 : _GEN_7339; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7670 = cnt[0] ? _GEN_7660 : _GEN_7340; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7671 = cnt[0] ? _GEN_7661 : _GEN_7341; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7672 = cnt[0] ? _GEN_7662 : _GEN_7342; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7673 = cnt[0] ? _GEN_7663 : _GEN_7343; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7674 = cnt[0] ? _GEN_7664 : _GEN_7344; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7675 = cnt[0] ? _GEN_7665 : _GEN_7345; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7676 = cnt[0] ? _GEN_7666 : _GEN_7346; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_7677 = cnt[0] ? _GEN_7667 : _GEN_7347; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7679 = _GEN_145 | _GEN_7669; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7680 = _GEN_146 | _GEN_7670; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7681 = _GEN_147 | _GEN_7671; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7682 = _GEN_148 | _GEN_7672; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_7683 = 2'h0 == opidx ? 5'h6 : _GEN_7673; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7684 = 2'h1 == opidx ? 5'h6 : _GEN_7674; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7685 = 2'h2 == opidx ? 5'h6 : _GEN_7675; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7686 = 2'h3 == opidx ? 5'h6 : _GEN_7676; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_7687 = _T_122 ? _cnt_T : _GEN_7677; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_7689 = cnt[1] ? _GEN_7679 : _GEN_7669; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7690 = cnt[1] ? _GEN_7680 : _GEN_7670; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7691 = cnt[1] ? _GEN_7681 : _GEN_7671; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7692 = cnt[1] ? _GEN_7682 : _GEN_7672; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7693 = cnt[1] ? _GEN_7683 : _GEN_7673; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7694 = cnt[1] ? _GEN_7684 : _GEN_7674; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7695 = cnt[1] ? _GEN_7685 : _GEN_7675; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7696 = cnt[1] ? _GEN_7686 : _GEN_7676; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_7697 = cnt[1] ? _GEN_7687 : _GEN_7677; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7699 = _GEN_145 | _GEN_7689; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7700 = _GEN_146 | _GEN_7690; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7701 = _GEN_147 | _GEN_7691; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7702 = _GEN_148 | _GEN_7692; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_7703 = 2'h0 == opidx ? 5'h7 : _GEN_7693; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7704 = 2'h1 == opidx ? 5'h7 : _GEN_7694; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7705 = 2'h2 == opidx ? 5'h7 : _GEN_7695; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7706 = 2'h3 == opidx ? 5'h7 : _GEN_7696; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_7707 = _T_122 ? _cnt_T : _GEN_7697; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_7709 = cnt[2] ? _GEN_7699 : _GEN_7689; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7710 = cnt[2] ? _GEN_7700 : _GEN_7690; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7711 = cnt[2] ? _GEN_7701 : _GEN_7691; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7712 = cnt[2] ? _GEN_7702 : _GEN_7692; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7713 = cnt[2] ? _GEN_7703 : _GEN_7693; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7714 = cnt[2] ? _GEN_7704 : _GEN_7694; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7715 = cnt[2] ? _GEN_7705 : _GEN_7695; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7716 = cnt[2] ? _GEN_7706 : _GEN_7696; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_7717 = cnt[2] ? _GEN_7707 : _GEN_7697; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7719 = _GEN_145 | _GEN_7709; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7720 = _GEN_146 | _GEN_7710; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7721 = _GEN_147 | _GEN_7711; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7722 = _GEN_148 | _GEN_7712; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_7723 = 2'h0 == opidx ? 5'h8 : _GEN_7713; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7724 = 2'h1 == opidx ? 5'h8 : _GEN_7714; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7725 = 2'h2 == opidx ? 5'h8 : _GEN_7715; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7726 = 2'h3 == opidx ? 5'h8 : _GEN_7716; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_7727 = _T_122 ? _cnt_T : _GEN_7717; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_7729 = cnt[3] ? _GEN_7719 : _GEN_7709; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7730 = cnt[3] ? _GEN_7720 : _GEN_7710; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7731 = cnt[3] ? _GEN_7721 : _GEN_7711; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7732 = cnt[3] ? _GEN_7722 : _GEN_7712; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7733 = cnt[3] ? _GEN_7723 : _GEN_7713; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7734 = cnt[3] ? _GEN_7724 : _GEN_7714; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7735 = cnt[3] ? _GEN_7725 : _GEN_7715; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7736 = cnt[3] ? _GEN_7726 : _GEN_7716; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_7737 = cnt[3] ? _GEN_7727 : _GEN_7717; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7739 = _GEN_145 | _GEN_7729; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7740 = _GEN_146 | _GEN_7730; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7741 = _GEN_147 | _GEN_7731; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7742 = _GEN_148 | _GEN_7732; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_7743 = 2'h0 == opidx ? 5'h9 : _GEN_7733; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7744 = 2'h1 == opidx ? 5'h9 : _GEN_7734; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7745 = 2'h2 == opidx ? 5'h9 : _GEN_7735; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7746 = 2'h3 == opidx ? 5'h9 : _GEN_7736; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_7747 = _T_122 ? _cnt_T : _GEN_7737; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_7749 = cnt[4] ? _GEN_7739 : _GEN_7729; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7750 = cnt[4] ? _GEN_7740 : _GEN_7730; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7751 = cnt[4] ? _GEN_7741 : _GEN_7731; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7752 = cnt[4] ? _GEN_7742 : _GEN_7732; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7753 = cnt[4] ? _GEN_7743 : _GEN_7733; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7754 = cnt[4] ? _GEN_7744 : _GEN_7734; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7755 = cnt[4] ? _GEN_7745 : _GEN_7735; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7756 = cnt[4] ? _GEN_7746 : _GEN_7736; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_7757 = cnt[4] ? _GEN_7747 : _GEN_7737; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7759 = _GEN_145 | _GEN_7749; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7760 = _GEN_146 | _GEN_7750; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7761 = _GEN_147 | _GEN_7751; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7762 = _GEN_148 | _GEN_7752; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_7763 = 2'h0 == opidx ? 5'ha : _GEN_7753; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7764 = 2'h1 == opidx ? 5'ha : _GEN_7754; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7765 = 2'h2 == opidx ? 5'ha : _GEN_7755; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7766 = 2'h3 == opidx ? 5'ha : _GEN_7756; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_7767 = _T_122 ? _cnt_T : _GEN_7757; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_7769 = cnt[5] ? _GEN_7759 : _GEN_7749; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7770 = cnt[5] ? _GEN_7760 : _GEN_7750; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7771 = cnt[5] ? _GEN_7761 : _GEN_7751; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7772 = cnt[5] ? _GEN_7762 : _GEN_7752; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7773 = cnt[5] ? _GEN_7763 : _GEN_7753; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7774 = cnt[5] ? _GEN_7764 : _GEN_7754; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7775 = cnt[5] ? _GEN_7765 : _GEN_7755; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7776 = cnt[5] ? _GEN_7766 : _GEN_7756; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_7777 = cnt[5] ? _GEN_7767 : _GEN_7757; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7779 = _GEN_145 | _GEN_7769; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7780 = _GEN_146 | _GEN_7770; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7781 = _GEN_147 | _GEN_7771; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7782 = _GEN_148 | _GEN_7772; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_7783 = 2'h0 == opidx ? 5'hb : _GEN_7773; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7784 = 2'h1 == opidx ? 5'hb : _GEN_7774; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7785 = 2'h2 == opidx ? 5'hb : _GEN_7775; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7786 = 2'h3 == opidx ? 5'hb : _GEN_7776; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_7787 = _T_122 ? _cnt_T : _GEN_7777; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_7789 = cnt[6] ? _GEN_7779 : _GEN_7769; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7790 = cnt[6] ? _GEN_7780 : _GEN_7770; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7791 = cnt[6] ? _GEN_7781 : _GEN_7771; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7792 = cnt[6] ? _GEN_7782 : _GEN_7772; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7793 = cnt[6] ? _GEN_7783 : _GEN_7773; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7794 = cnt[6] ? _GEN_7784 : _GEN_7774; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7795 = cnt[6] ? _GEN_7785 : _GEN_7775; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7796 = cnt[6] ? _GEN_7786 : _GEN_7776; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_7797 = cnt[6] ? _GEN_7787 : _GEN_7777; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7799 = _GEN_145 | _GEN_7789; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7800 = _GEN_146 | _GEN_7790; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7801 = _GEN_147 | _GEN_7791; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7802 = _GEN_148 | _GEN_7792; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_7803 = 2'h0 == opidx ? 5'hc : _GEN_7793; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7804 = 2'h1 == opidx ? 5'hc : _GEN_7794; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7805 = 2'h2 == opidx ? 5'hc : _GEN_7795; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7806 = 2'h3 == opidx ? 5'hc : _GEN_7796; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_7807 = _T_122 ? _cnt_T : _GEN_7797; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_7809 = cnt[7] ? _GEN_7799 : _GEN_7789; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7810 = cnt[7] ? _GEN_7800 : _GEN_7790; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7811 = cnt[7] ? _GEN_7801 : _GEN_7791; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7812 = cnt[7] ? _GEN_7802 : _GEN_7792; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7813 = cnt[7] ? _GEN_7803 : _GEN_7793; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7814 = cnt[7] ? _GEN_7804 : _GEN_7794; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7815 = cnt[7] ? _GEN_7805 : _GEN_7795; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7816 = cnt[7] ? _GEN_7806 : _GEN_7796; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_7817 = cnt[7] ? _GEN_7807 : _GEN_7797; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7819 = _GEN_145 | _GEN_7809; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7820 = _GEN_146 | _GEN_7810; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7821 = _GEN_147 | _GEN_7811; // @[NulCtrlMP.scala 351:{27,27}]
  wire  _GEN_7822 = _GEN_148 | _GEN_7812; // @[NulCtrlMP.scala 351:{27,27}]
  wire [4:0] _GEN_7823 = 2'h0 == opidx ? 5'hd : _GEN_7813; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7824 = 2'h1 == opidx ? 5'hd : _GEN_7814; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7825 = 2'h2 == opidx ? 5'hd : _GEN_7815; // @[NulCtrlMP.scala 352:{28,28}]
  wire [4:0] _GEN_7826 = 2'h3 == opidx ? 5'hd : _GEN_7816; // @[NulCtrlMP.scala 352:{28,28}]
  wire [128:0] _GEN_7827 = _T_122 ? _cnt_T : _GEN_7817; // @[NulCtrlMP.scala 353:36 354:17]
  wire  _GEN_7829 = cnt[8] ? _GEN_7819 : _GEN_7809; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7830 = cnt[8] ? _GEN_7820 : _GEN_7810; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7831 = cnt[8] ? _GEN_7821 : _GEN_7811; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7832 = cnt[8] ? _GEN_7822 : _GEN_7812; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7833 = cnt[8] ? _GEN_7823 : _GEN_7813; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7834 = cnt[8] ? _GEN_7824 : _GEN_7814; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7835 = cnt[8] ? _GEN_7825 : _GEN_7815; // @[NulCtrlMP.scala 408:32]
  wire [4:0] _GEN_7836 = cnt[8] ? _GEN_7826 : _GEN_7816; // @[NulCtrlMP.scala 408:32]
  wire [128:0] _GEN_7837 = cnt[8] ? _GEN_7827 : _GEN_7817; // @[NulCtrlMP.scala 408:32]
  wire  _GEN_7839 = _GEN_145 | _GEN_7359; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7840 = _GEN_146 | _GEN_7360; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7841 = _GEN_147 | _GEN_7361; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7842 = _GEN_148 | _GEN_7362; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7843 = 2'h0 == opidx ? 5'h5 : _GEN_7833; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7844 = 2'h1 == opidx ? 5'h5 : _GEN_7834; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7845 = 2'h2 == opidx ? 5'h5 : _GEN_7835; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7846 = 2'h3 == opidx ? 5'h5 : _GEN_7836; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7847 = 2'h0 == opidx ? _T_464 : _GEN_7363; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7848 = 2'h1 == opidx ? _T_464 : _GEN_7364; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7849 = 2'h2 == opidx ? _T_464 : _GEN_7365; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7850 = 2'h3 == opidx ? _T_464 : _GEN_7366; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7851 = ~_GEN_1128 ? _cnt_T : _GEN_7837; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7852 = cnt[9] ? _GEN_7839 : _GEN_7359; // @[NulCtrlMP.scala 895:22]
  wire  _GEN_7853 = cnt[9] ? _GEN_7840 : _GEN_7360; // @[NulCtrlMP.scala 895:22]
  wire  _GEN_7854 = cnt[9] ? _GEN_7841 : _GEN_7361; // @[NulCtrlMP.scala 895:22]
  wire  _GEN_7855 = cnt[9] ? _GEN_7842 : _GEN_7362; // @[NulCtrlMP.scala 895:22]
  wire [4:0] _GEN_7856 = cnt[9] ? _GEN_7843 : _GEN_7833; // @[NulCtrlMP.scala 895:22]
  wire [4:0] _GEN_7857 = cnt[9] ? _GEN_7844 : _GEN_7834; // @[NulCtrlMP.scala 895:22]
  wire [4:0] _GEN_7858 = cnt[9] ? _GEN_7845 : _GEN_7835; // @[NulCtrlMP.scala 895:22]
  wire [4:0] _GEN_7859 = cnt[9] ? _GEN_7846 : _GEN_7836; // @[NulCtrlMP.scala 895:22]
  wire [63:0] _GEN_7860 = cnt[9] ? _GEN_7847 : _GEN_7363; // @[NulCtrlMP.scala 895:22]
  wire [63:0] _GEN_7861 = cnt[9] ? _GEN_7848 : _GEN_7364; // @[NulCtrlMP.scala 895:22]
  wire [63:0] _GEN_7862 = cnt[9] ? _GEN_7849 : _GEN_7365; // @[NulCtrlMP.scala 895:22]
  wire [63:0] _GEN_7863 = cnt[9] ? _GEN_7850 : _GEN_7366; // @[NulCtrlMP.scala 895:22]
  wire [128:0] _GEN_7864 = cnt[9] ? _GEN_7851 : _GEN_7837; // @[NulCtrlMP.scala 895:22]
  wire [128:0] _GEN_7865 = pgbuf_uart_pos >= _pgbuf_cpu_pos_T_1 ? _cnt_T : _GEN_7864; // @[NulCtrlMP.scala 897:58 898:21]
  wire [128:0] _GEN_7866 = cnt[10] ? _GEN_7865 : _GEN_7864; // @[NulCtrlMP.scala 896:23]
  wire  _GEN_7867 = _GEN_145 | _GEN_7852; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7868 = _GEN_146 | _GEN_7853; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7869 = _GEN_147 | _GEN_7854; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7870 = _GEN_148 | _GEN_7855; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7871 = 2'h0 == opidx ? 5'h6 : _GEN_7856; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7872 = 2'h1 == opidx ? 5'h6 : _GEN_7857; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7873 = 2'h2 == opidx ? 5'h6 : _GEN_7858; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7874 = 2'h3 == opidx ? 5'h6 : _GEN_7859; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7880 = 6'h1 == _T_479[5:0] ? pgbuf_div8_1 : pgbuf_div8_0; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7881 = 6'h2 == _T_479[5:0] ? pgbuf_div8_2 : _GEN_7880; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7882 = 6'h3 == _T_479[5:0] ? pgbuf_div8_3 : _GEN_7881; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7883 = 6'h4 == _T_479[5:0] ? pgbuf_div8_4 : _GEN_7882; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7884 = 6'h5 == _T_479[5:0] ? pgbuf_div8_5 : _GEN_7883; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7885 = 6'h6 == _T_479[5:0] ? pgbuf_div8_6 : _GEN_7884; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7886 = 6'h7 == _T_479[5:0] ? pgbuf_div8_7 : _GEN_7885; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7887 = 6'h8 == _T_479[5:0] ? pgbuf_div8_8 : _GEN_7886; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7888 = 6'h9 == _T_479[5:0] ? pgbuf_div8_9 : _GEN_7887; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7889 = 6'ha == _T_479[5:0] ? pgbuf_div8_10 : _GEN_7888; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7890 = 6'hb == _T_479[5:0] ? pgbuf_div8_11 : _GEN_7889; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7891 = 6'hc == _T_479[5:0] ? pgbuf_div8_12 : _GEN_7890; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7892 = 6'hd == _T_479[5:0] ? pgbuf_div8_13 : _GEN_7891; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7893 = 6'he == _T_479[5:0] ? pgbuf_div8_14 : _GEN_7892; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7894 = 6'hf == _T_479[5:0] ? pgbuf_div8_15 : _GEN_7893; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7895 = 6'h10 == _T_479[5:0] ? pgbuf_div8_16 : _GEN_7894; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7896 = 6'h11 == _T_479[5:0] ? pgbuf_div8_17 : _GEN_7895; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7897 = 6'h12 == _T_479[5:0] ? pgbuf_div8_18 : _GEN_7896; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7898 = 6'h13 == _T_479[5:0] ? pgbuf_div8_19 : _GEN_7897; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7899 = 6'h14 == _T_479[5:0] ? pgbuf_div8_20 : _GEN_7898; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7900 = 6'h15 == _T_479[5:0] ? pgbuf_div8_21 : _GEN_7899; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7901 = 6'h16 == _T_479[5:0] ? pgbuf_div8_22 : _GEN_7900; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7902 = 6'h17 == _T_479[5:0] ? pgbuf_div8_23 : _GEN_7901; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7903 = 6'h18 == _T_479[5:0] ? pgbuf_div8_24 : _GEN_7902; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7904 = 6'h19 == _T_479[5:0] ? pgbuf_div8_25 : _GEN_7903; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7905 = 6'h1a == _T_479[5:0] ? pgbuf_div8_26 : _GEN_7904; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7906 = 6'h1b == _T_479[5:0] ? pgbuf_div8_27 : _GEN_7905; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7907 = 6'h1c == _T_479[5:0] ? pgbuf_div8_28 : _GEN_7906; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7908 = 6'h1d == _T_479[5:0] ? pgbuf_div8_29 : _GEN_7907; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7909 = 6'h1e == _T_479[5:0] ? pgbuf_div8_30 : _GEN_7908; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7910 = 6'h1f == _T_479[5:0] ? pgbuf_div8_31 : _GEN_7909; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7911 = 6'h20 == _T_479[5:0] ? pgbuf_div8_32 : _GEN_7910; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7912 = 6'h21 == _T_479[5:0] ? pgbuf_div8_33 : _GEN_7911; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7913 = 6'h22 == _T_479[5:0] ? pgbuf_div8_34 : _GEN_7912; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7914 = 6'h23 == _T_479[5:0] ? pgbuf_div8_35 : _GEN_7913; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7915 = 6'h24 == _T_479[5:0] ? pgbuf_div8_36 : _GEN_7914; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7916 = 6'h25 == _T_479[5:0] ? pgbuf_div8_37 : _GEN_7915; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7917 = 6'h26 == _T_479[5:0] ? pgbuf_div8_38 : _GEN_7916; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7918 = 6'h27 == _T_479[5:0] ? pgbuf_div8_39 : _GEN_7917; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7919 = 6'h28 == _T_479[5:0] ? pgbuf_div8_40 : _GEN_7918; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7920 = 6'h29 == _T_479[5:0] ? pgbuf_div8_41 : _GEN_7919; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7921 = 6'h2a == _T_479[5:0] ? pgbuf_div8_42 : _GEN_7920; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7922 = 6'h2b == _T_479[5:0] ? pgbuf_div8_43 : _GEN_7921; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7923 = 6'h2c == _T_479[5:0] ? pgbuf_div8_44 : _GEN_7922; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7924 = 6'h2d == _T_479[5:0] ? pgbuf_div8_45 : _GEN_7923; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7925 = 6'h2e == _T_479[5:0] ? pgbuf_div8_46 : _GEN_7924; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7926 = 6'h2f == _T_479[5:0] ? pgbuf_div8_47 : _GEN_7925; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7927 = 6'h30 == _T_479[5:0] ? pgbuf_div8_48 : _GEN_7926; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7928 = 6'h31 == _T_479[5:0] ? pgbuf_div8_49 : _GEN_7927; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7929 = 6'h32 == _T_479[5:0] ? pgbuf_div8_50 : _GEN_7928; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7930 = 6'h33 == _T_479[5:0] ? pgbuf_div8_51 : _GEN_7929; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7931 = 6'h34 == _T_479[5:0] ? pgbuf_div8_52 : _GEN_7930; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7932 = 6'h35 == _T_479[5:0] ? pgbuf_div8_53 : _GEN_7931; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7933 = 6'h36 == _T_479[5:0] ? pgbuf_div8_54 : _GEN_7932; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7934 = 6'h37 == _T_479[5:0] ? pgbuf_div8_55 : _GEN_7933; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7935 = 6'h38 == _T_479[5:0] ? pgbuf_div8_56 : _GEN_7934; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7936 = 6'h39 == _T_479[5:0] ? pgbuf_div8_57 : _GEN_7935; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7937 = 6'h3a == _T_479[5:0] ? pgbuf_div8_58 : _GEN_7936; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7938 = 6'h3b == _T_479[5:0] ? pgbuf_div8_59 : _GEN_7937; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7939 = 6'h3c == _T_479[5:0] ? pgbuf_div8_60 : _GEN_7938; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7940 = 6'h3d == _T_479[5:0] ? pgbuf_div8_61 : _GEN_7939; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7941 = 6'h3e == _T_479[5:0] ? pgbuf_div8_62 : _GEN_7940; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7942 = 6'h3f == _T_479[5:0] ? pgbuf_div8_63 : _GEN_7941; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7875 = 2'h0 == opidx ? _GEN_7942 : _GEN_7860; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7876 = 2'h1 == opidx ? _GEN_7942 : _GEN_7861; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7877 = 2'h2 == opidx ? _GEN_7942 : _GEN_7862; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7878 = 2'h3 == opidx ? _GEN_7942 : _GEN_7863; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_7943 = ~_GEN_1128 ? _cnt_T : _GEN_7866; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_7944 = cnt[11] ? _GEN_7867 : _GEN_7852; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_7945 = cnt[11] ? _GEN_7868 : _GEN_7853; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_7946 = cnt[11] ? _GEN_7869 : _GEN_7854; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_7947 = cnt[11] ? _GEN_7870 : _GEN_7855; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_7948 = cnt[11] ? _GEN_7871 : _GEN_7856; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_7949 = cnt[11] ? _GEN_7872 : _GEN_7857; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_7950 = cnt[11] ? _GEN_7873 : _GEN_7858; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_7951 = cnt[11] ? _GEN_7874 : _GEN_7859; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_7952 = cnt[11] ? _GEN_7875 : _GEN_7860; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_7953 = cnt[11] ? _GEN_7876 : _GEN_7861; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_7954 = cnt[11] ? _GEN_7877 : _GEN_7862; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_7955 = cnt[11] ? _GEN_7878 : _GEN_7863; // @[NulCtrlMP.scala 902:29]
  wire [128:0] _GEN_7956 = cnt[11] ? _GEN_7943 : _GEN_7866; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_7957 = _GEN_145 | _GEN_7944; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7958 = _GEN_146 | _GEN_7945; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7959 = _GEN_147 | _GEN_7946; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_7960 = _GEN_148 | _GEN_7947; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_7961 = 2'h0 == opidx ? 5'h7 : _GEN_7948; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7962 = 2'h1 == opidx ? 5'h7 : _GEN_7949; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7963 = 2'h2 == opidx ? 5'h7 : _GEN_7950; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_7964 = 2'h3 == opidx ? 5'h7 : _GEN_7951; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_7970 = 6'h1 == _T_486[5:0] ? pgbuf_div8_1 : pgbuf_div8_0; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7971 = 6'h2 == _T_486[5:0] ? pgbuf_div8_2 : _GEN_7970; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7972 = 6'h3 == _T_486[5:0] ? pgbuf_div8_3 : _GEN_7971; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7973 = 6'h4 == _T_486[5:0] ? pgbuf_div8_4 : _GEN_7972; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7974 = 6'h5 == _T_486[5:0] ? pgbuf_div8_5 : _GEN_7973; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7975 = 6'h6 == _T_486[5:0] ? pgbuf_div8_6 : _GEN_7974; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7976 = 6'h7 == _T_486[5:0] ? pgbuf_div8_7 : _GEN_7975; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7977 = 6'h8 == _T_486[5:0] ? pgbuf_div8_8 : _GEN_7976; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7978 = 6'h9 == _T_486[5:0] ? pgbuf_div8_9 : _GEN_7977; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7979 = 6'ha == _T_486[5:0] ? pgbuf_div8_10 : _GEN_7978; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7980 = 6'hb == _T_486[5:0] ? pgbuf_div8_11 : _GEN_7979; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7981 = 6'hc == _T_486[5:0] ? pgbuf_div8_12 : _GEN_7980; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7982 = 6'hd == _T_486[5:0] ? pgbuf_div8_13 : _GEN_7981; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7983 = 6'he == _T_486[5:0] ? pgbuf_div8_14 : _GEN_7982; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7984 = 6'hf == _T_486[5:0] ? pgbuf_div8_15 : _GEN_7983; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7985 = 6'h10 == _T_486[5:0] ? pgbuf_div8_16 : _GEN_7984; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7986 = 6'h11 == _T_486[5:0] ? pgbuf_div8_17 : _GEN_7985; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7987 = 6'h12 == _T_486[5:0] ? pgbuf_div8_18 : _GEN_7986; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7988 = 6'h13 == _T_486[5:0] ? pgbuf_div8_19 : _GEN_7987; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7989 = 6'h14 == _T_486[5:0] ? pgbuf_div8_20 : _GEN_7988; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7990 = 6'h15 == _T_486[5:0] ? pgbuf_div8_21 : _GEN_7989; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7991 = 6'h16 == _T_486[5:0] ? pgbuf_div8_22 : _GEN_7990; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7992 = 6'h17 == _T_486[5:0] ? pgbuf_div8_23 : _GEN_7991; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7993 = 6'h18 == _T_486[5:0] ? pgbuf_div8_24 : _GEN_7992; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7994 = 6'h19 == _T_486[5:0] ? pgbuf_div8_25 : _GEN_7993; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7995 = 6'h1a == _T_486[5:0] ? pgbuf_div8_26 : _GEN_7994; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7996 = 6'h1b == _T_486[5:0] ? pgbuf_div8_27 : _GEN_7995; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7997 = 6'h1c == _T_486[5:0] ? pgbuf_div8_28 : _GEN_7996; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7998 = 6'h1d == _T_486[5:0] ? pgbuf_div8_29 : _GEN_7997; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7999 = 6'h1e == _T_486[5:0] ? pgbuf_div8_30 : _GEN_7998; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8000 = 6'h1f == _T_486[5:0] ? pgbuf_div8_31 : _GEN_7999; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8001 = 6'h20 == _T_486[5:0] ? pgbuf_div8_32 : _GEN_8000; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8002 = 6'h21 == _T_486[5:0] ? pgbuf_div8_33 : _GEN_8001; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8003 = 6'h22 == _T_486[5:0] ? pgbuf_div8_34 : _GEN_8002; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8004 = 6'h23 == _T_486[5:0] ? pgbuf_div8_35 : _GEN_8003; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8005 = 6'h24 == _T_486[5:0] ? pgbuf_div8_36 : _GEN_8004; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8006 = 6'h25 == _T_486[5:0] ? pgbuf_div8_37 : _GEN_8005; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8007 = 6'h26 == _T_486[5:0] ? pgbuf_div8_38 : _GEN_8006; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8008 = 6'h27 == _T_486[5:0] ? pgbuf_div8_39 : _GEN_8007; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8009 = 6'h28 == _T_486[5:0] ? pgbuf_div8_40 : _GEN_8008; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8010 = 6'h29 == _T_486[5:0] ? pgbuf_div8_41 : _GEN_8009; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8011 = 6'h2a == _T_486[5:0] ? pgbuf_div8_42 : _GEN_8010; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8012 = 6'h2b == _T_486[5:0] ? pgbuf_div8_43 : _GEN_8011; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8013 = 6'h2c == _T_486[5:0] ? pgbuf_div8_44 : _GEN_8012; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8014 = 6'h2d == _T_486[5:0] ? pgbuf_div8_45 : _GEN_8013; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8015 = 6'h2e == _T_486[5:0] ? pgbuf_div8_46 : _GEN_8014; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8016 = 6'h2f == _T_486[5:0] ? pgbuf_div8_47 : _GEN_8015; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8017 = 6'h30 == _T_486[5:0] ? pgbuf_div8_48 : _GEN_8016; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8018 = 6'h31 == _T_486[5:0] ? pgbuf_div8_49 : _GEN_8017; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8019 = 6'h32 == _T_486[5:0] ? pgbuf_div8_50 : _GEN_8018; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8020 = 6'h33 == _T_486[5:0] ? pgbuf_div8_51 : _GEN_8019; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8021 = 6'h34 == _T_486[5:0] ? pgbuf_div8_52 : _GEN_8020; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8022 = 6'h35 == _T_486[5:0] ? pgbuf_div8_53 : _GEN_8021; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8023 = 6'h36 == _T_486[5:0] ? pgbuf_div8_54 : _GEN_8022; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8024 = 6'h37 == _T_486[5:0] ? pgbuf_div8_55 : _GEN_8023; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8025 = 6'h38 == _T_486[5:0] ? pgbuf_div8_56 : _GEN_8024; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8026 = 6'h39 == _T_486[5:0] ? pgbuf_div8_57 : _GEN_8025; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8027 = 6'h3a == _T_486[5:0] ? pgbuf_div8_58 : _GEN_8026; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8028 = 6'h3b == _T_486[5:0] ? pgbuf_div8_59 : _GEN_8027; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8029 = 6'h3c == _T_486[5:0] ? pgbuf_div8_60 : _GEN_8028; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8030 = 6'h3d == _T_486[5:0] ? pgbuf_div8_61 : _GEN_8029; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8031 = 6'h3e == _T_486[5:0] ? pgbuf_div8_62 : _GEN_8030; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8032 = 6'h3f == _T_486[5:0] ? pgbuf_div8_63 : _GEN_8031; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7965 = 2'h0 == opidx ? _GEN_8032 : _GEN_7952; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7966 = 2'h1 == opidx ? _GEN_8032 : _GEN_7953; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7967 = 2'h2 == opidx ? _GEN_8032 : _GEN_7954; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_7968 = 2'h3 == opidx ? _GEN_8032 : _GEN_7955; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8033 = ~_GEN_1128 ? _cnt_T : _GEN_7956; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8034 = cnt[12] ? _GEN_7957 : _GEN_7944; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8035 = cnt[12] ? _GEN_7958 : _GEN_7945; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8036 = cnt[12] ? _GEN_7959 : _GEN_7946; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8037 = cnt[12] ? _GEN_7960 : _GEN_7947; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8038 = cnt[12] ? _GEN_7961 : _GEN_7948; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8039 = cnt[12] ? _GEN_7962 : _GEN_7949; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8040 = cnt[12] ? _GEN_7963 : _GEN_7950; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8041 = cnt[12] ? _GEN_7964 : _GEN_7951; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8042 = cnt[12] ? _GEN_7965 : _GEN_7952; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8043 = cnt[12] ? _GEN_7966 : _GEN_7953; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8044 = cnt[12] ? _GEN_7967 : _GEN_7954; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8045 = cnt[12] ? _GEN_7968 : _GEN_7955; // @[NulCtrlMP.scala 902:29]
  wire [128:0] _GEN_8046 = cnt[12] ? _GEN_8033 : _GEN_7956; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8047 = _GEN_145 | _GEN_8034; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8048 = _GEN_146 | _GEN_8035; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8049 = _GEN_147 | _GEN_8036; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8050 = _GEN_148 | _GEN_8037; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8051 = 2'h0 == opidx ? 5'h8 : _GEN_8038; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8052 = 2'h1 == opidx ? 5'h8 : _GEN_8039; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8053 = 2'h2 == opidx ? 5'h8 : _GEN_8040; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8054 = 2'h3 == opidx ? 5'h8 : _GEN_8041; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8060 = 6'h1 == _T_492[5:0] ? pgbuf_div8_1 : pgbuf_div8_0; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8061 = 6'h2 == _T_492[5:0] ? pgbuf_div8_2 : _GEN_8060; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8062 = 6'h3 == _T_492[5:0] ? pgbuf_div8_3 : _GEN_8061; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8063 = 6'h4 == _T_492[5:0] ? pgbuf_div8_4 : _GEN_8062; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8064 = 6'h5 == _T_492[5:0] ? pgbuf_div8_5 : _GEN_8063; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8065 = 6'h6 == _T_492[5:0] ? pgbuf_div8_6 : _GEN_8064; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8066 = 6'h7 == _T_492[5:0] ? pgbuf_div8_7 : _GEN_8065; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8067 = 6'h8 == _T_492[5:0] ? pgbuf_div8_8 : _GEN_8066; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8068 = 6'h9 == _T_492[5:0] ? pgbuf_div8_9 : _GEN_8067; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8069 = 6'ha == _T_492[5:0] ? pgbuf_div8_10 : _GEN_8068; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8070 = 6'hb == _T_492[5:0] ? pgbuf_div8_11 : _GEN_8069; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8071 = 6'hc == _T_492[5:0] ? pgbuf_div8_12 : _GEN_8070; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8072 = 6'hd == _T_492[5:0] ? pgbuf_div8_13 : _GEN_8071; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8073 = 6'he == _T_492[5:0] ? pgbuf_div8_14 : _GEN_8072; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8074 = 6'hf == _T_492[5:0] ? pgbuf_div8_15 : _GEN_8073; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8075 = 6'h10 == _T_492[5:0] ? pgbuf_div8_16 : _GEN_8074; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8076 = 6'h11 == _T_492[5:0] ? pgbuf_div8_17 : _GEN_8075; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8077 = 6'h12 == _T_492[5:0] ? pgbuf_div8_18 : _GEN_8076; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8078 = 6'h13 == _T_492[5:0] ? pgbuf_div8_19 : _GEN_8077; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8079 = 6'h14 == _T_492[5:0] ? pgbuf_div8_20 : _GEN_8078; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8080 = 6'h15 == _T_492[5:0] ? pgbuf_div8_21 : _GEN_8079; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8081 = 6'h16 == _T_492[5:0] ? pgbuf_div8_22 : _GEN_8080; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8082 = 6'h17 == _T_492[5:0] ? pgbuf_div8_23 : _GEN_8081; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8083 = 6'h18 == _T_492[5:0] ? pgbuf_div8_24 : _GEN_8082; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8084 = 6'h19 == _T_492[5:0] ? pgbuf_div8_25 : _GEN_8083; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8085 = 6'h1a == _T_492[5:0] ? pgbuf_div8_26 : _GEN_8084; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8086 = 6'h1b == _T_492[5:0] ? pgbuf_div8_27 : _GEN_8085; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8087 = 6'h1c == _T_492[5:0] ? pgbuf_div8_28 : _GEN_8086; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8088 = 6'h1d == _T_492[5:0] ? pgbuf_div8_29 : _GEN_8087; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8089 = 6'h1e == _T_492[5:0] ? pgbuf_div8_30 : _GEN_8088; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8090 = 6'h1f == _T_492[5:0] ? pgbuf_div8_31 : _GEN_8089; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8091 = 6'h20 == _T_492[5:0] ? pgbuf_div8_32 : _GEN_8090; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8092 = 6'h21 == _T_492[5:0] ? pgbuf_div8_33 : _GEN_8091; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8093 = 6'h22 == _T_492[5:0] ? pgbuf_div8_34 : _GEN_8092; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8094 = 6'h23 == _T_492[5:0] ? pgbuf_div8_35 : _GEN_8093; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8095 = 6'h24 == _T_492[5:0] ? pgbuf_div8_36 : _GEN_8094; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8096 = 6'h25 == _T_492[5:0] ? pgbuf_div8_37 : _GEN_8095; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8097 = 6'h26 == _T_492[5:0] ? pgbuf_div8_38 : _GEN_8096; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8098 = 6'h27 == _T_492[5:0] ? pgbuf_div8_39 : _GEN_8097; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8099 = 6'h28 == _T_492[5:0] ? pgbuf_div8_40 : _GEN_8098; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8100 = 6'h29 == _T_492[5:0] ? pgbuf_div8_41 : _GEN_8099; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8101 = 6'h2a == _T_492[5:0] ? pgbuf_div8_42 : _GEN_8100; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8102 = 6'h2b == _T_492[5:0] ? pgbuf_div8_43 : _GEN_8101; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8103 = 6'h2c == _T_492[5:0] ? pgbuf_div8_44 : _GEN_8102; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8104 = 6'h2d == _T_492[5:0] ? pgbuf_div8_45 : _GEN_8103; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8105 = 6'h2e == _T_492[5:0] ? pgbuf_div8_46 : _GEN_8104; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8106 = 6'h2f == _T_492[5:0] ? pgbuf_div8_47 : _GEN_8105; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8107 = 6'h30 == _T_492[5:0] ? pgbuf_div8_48 : _GEN_8106; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8108 = 6'h31 == _T_492[5:0] ? pgbuf_div8_49 : _GEN_8107; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8109 = 6'h32 == _T_492[5:0] ? pgbuf_div8_50 : _GEN_8108; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8110 = 6'h33 == _T_492[5:0] ? pgbuf_div8_51 : _GEN_8109; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8111 = 6'h34 == _T_492[5:0] ? pgbuf_div8_52 : _GEN_8110; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8112 = 6'h35 == _T_492[5:0] ? pgbuf_div8_53 : _GEN_8111; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8113 = 6'h36 == _T_492[5:0] ? pgbuf_div8_54 : _GEN_8112; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8114 = 6'h37 == _T_492[5:0] ? pgbuf_div8_55 : _GEN_8113; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8115 = 6'h38 == _T_492[5:0] ? pgbuf_div8_56 : _GEN_8114; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8116 = 6'h39 == _T_492[5:0] ? pgbuf_div8_57 : _GEN_8115; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8117 = 6'h3a == _T_492[5:0] ? pgbuf_div8_58 : _GEN_8116; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8118 = 6'h3b == _T_492[5:0] ? pgbuf_div8_59 : _GEN_8117; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8119 = 6'h3c == _T_492[5:0] ? pgbuf_div8_60 : _GEN_8118; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8120 = 6'h3d == _T_492[5:0] ? pgbuf_div8_61 : _GEN_8119; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8121 = 6'h3e == _T_492[5:0] ? pgbuf_div8_62 : _GEN_8120; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8122 = 6'h3f == _T_492[5:0] ? pgbuf_div8_63 : _GEN_8121; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8055 = 2'h0 == opidx ? _GEN_8122 : _GEN_8042; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8056 = 2'h1 == opidx ? _GEN_8122 : _GEN_8043; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8057 = 2'h2 == opidx ? _GEN_8122 : _GEN_8044; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8058 = 2'h3 == opidx ? _GEN_8122 : _GEN_8045; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8123 = ~_GEN_1128 ? _cnt_T : _GEN_8046; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8124 = cnt[13] ? _GEN_8047 : _GEN_8034; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8125 = cnt[13] ? _GEN_8048 : _GEN_8035; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8126 = cnt[13] ? _GEN_8049 : _GEN_8036; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8127 = cnt[13] ? _GEN_8050 : _GEN_8037; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8128 = cnt[13] ? _GEN_8051 : _GEN_8038; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8129 = cnt[13] ? _GEN_8052 : _GEN_8039; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8130 = cnt[13] ? _GEN_8053 : _GEN_8040; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8131 = cnt[13] ? _GEN_8054 : _GEN_8041; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8132 = cnt[13] ? _GEN_8055 : _GEN_8042; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8133 = cnt[13] ? _GEN_8056 : _GEN_8043; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8134 = cnt[13] ? _GEN_8057 : _GEN_8044; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8135 = cnt[13] ? _GEN_8058 : _GEN_8045; // @[NulCtrlMP.scala 902:29]
  wire [128:0] _GEN_8136 = cnt[13] ? _GEN_8123 : _GEN_8046; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8137 = _GEN_145 | _GEN_8124; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8138 = _GEN_146 | _GEN_8125; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8139 = _GEN_147 | _GEN_8126; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8140 = _GEN_148 | _GEN_8127; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8141 = 2'h0 == opidx ? 5'h9 : _GEN_8128; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8142 = 2'h1 == opidx ? 5'h9 : _GEN_8129; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8143 = 2'h2 == opidx ? 5'h9 : _GEN_8130; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8144 = 2'h3 == opidx ? 5'h9 : _GEN_8131; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8150 = 6'h1 == _T_498[5:0] ? pgbuf_div8_1 : pgbuf_div8_0; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8151 = 6'h2 == _T_498[5:0] ? pgbuf_div8_2 : _GEN_8150; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8152 = 6'h3 == _T_498[5:0] ? pgbuf_div8_3 : _GEN_8151; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8153 = 6'h4 == _T_498[5:0] ? pgbuf_div8_4 : _GEN_8152; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8154 = 6'h5 == _T_498[5:0] ? pgbuf_div8_5 : _GEN_8153; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8155 = 6'h6 == _T_498[5:0] ? pgbuf_div8_6 : _GEN_8154; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8156 = 6'h7 == _T_498[5:0] ? pgbuf_div8_7 : _GEN_8155; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8157 = 6'h8 == _T_498[5:0] ? pgbuf_div8_8 : _GEN_8156; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8158 = 6'h9 == _T_498[5:0] ? pgbuf_div8_9 : _GEN_8157; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8159 = 6'ha == _T_498[5:0] ? pgbuf_div8_10 : _GEN_8158; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8160 = 6'hb == _T_498[5:0] ? pgbuf_div8_11 : _GEN_8159; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8161 = 6'hc == _T_498[5:0] ? pgbuf_div8_12 : _GEN_8160; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8162 = 6'hd == _T_498[5:0] ? pgbuf_div8_13 : _GEN_8161; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8163 = 6'he == _T_498[5:0] ? pgbuf_div8_14 : _GEN_8162; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8164 = 6'hf == _T_498[5:0] ? pgbuf_div8_15 : _GEN_8163; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8165 = 6'h10 == _T_498[5:0] ? pgbuf_div8_16 : _GEN_8164; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8166 = 6'h11 == _T_498[5:0] ? pgbuf_div8_17 : _GEN_8165; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8167 = 6'h12 == _T_498[5:0] ? pgbuf_div8_18 : _GEN_8166; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8168 = 6'h13 == _T_498[5:0] ? pgbuf_div8_19 : _GEN_8167; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8169 = 6'h14 == _T_498[5:0] ? pgbuf_div8_20 : _GEN_8168; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8170 = 6'h15 == _T_498[5:0] ? pgbuf_div8_21 : _GEN_8169; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8171 = 6'h16 == _T_498[5:0] ? pgbuf_div8_22 : _GEN_8170; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8172 = 6'h17 == _T_498[5:0] ? pgbuf_div8_23 : _GEN_8171; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8173 = 6'h18 == _T_498[5:0] ? pgbuf_div8_24 : _GEN_8172; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8174 = 6'h19 == _T_498[5:0] ? pgbuf_div8_25 : _GEN_8173; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8175 = 6'h1a == _T_498[5:0] ? pgbuf_div8_26 : _GEN_8174; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8176 = 6'h1b == _T_498[5:0] ? pgbuf_div8_27 : _GEN_8175; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8177 = 6'h1c == _T_498[5:0] ? pgbuf_div8_28 : _GEN_8176; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8178 = 6'h1d == _T_498[5:0] ? pgbuf_div8_29 : _GEN_8177; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8179 = 6'h1e == _T_498[5:0] ? pgbuf_div8_30 : _GEN_8178; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8180 = 6'h1f == _T_498[5:0] ? pgbuf_div8_31 : _GEN_8179; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8181 = 6'h20 == _T_498[5:0] ? pgbuf_div8_32 : _GEN_8180; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8182 = 6'h21 == _T_498[5:0] ? pgbuf_div8_33 : _GEN_8181; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8183 = 6'h22 == _T_498[5:0] ? pgbuf_div8_34 : _GEN_8182; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8184 = 6'h23 == _T_498[5:0] ? pgbuf_div8_35 : _GEN_8183; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8185 = 6'h24 == _T_498[5:0] ? pgbuf_div8_36 : _GEN_8184; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8186 = 6'h25 == _T_498[5:0] ? pgbuf_div8_37 : _GEN_8185; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8187 = 6'h26 == _T_498[5:0] ? pgbuf_div8_38 : _GEN_8186; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8188 = 6'h27 == _T_498[5:0] ? pgbuf_div8_39 : _GEN_8187; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8189 = 6'h28 == _T_498[5:0] ? pgbuf_div8_40 : _GEN_8188; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8190 = 6'h29 == _T_498[5:0] ? pgbuf_div8_41 : _GEN_8189; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8191 = 6'h2a == _T_498[5:0] ? pgbuf_div8_42 : _GEN_8190; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8192 = 6'h2b == _T_498[5:0] ? pgbuf_div8_43 : _GEN_8191; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8193 = 6'h2c == _T_498[5:0] ? pgbuf_div8_44 : _GEN_8192; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8194 = 6'h2d == _T_498[5:0] ? pgbuf_div8_45 : _GEN_8193; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8195 = 6'h2e == _T_498[5:0] ? pgbuf_div8_46 : _GEN_8194; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8196 = 6'h2f == _T_498[5:0] ? pgbuf_div8_47 : _GEN_8195; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8197 = 6'h30 == _T_498[5:0] ? pgbuf_div8_48 : _GEN_8196; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8198 = 6'h31 == _T_498[5:0] ? pgbuf_div8_49 : _GEN_8197; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8199 = 6'h32 == _T_498[5:0] ? pgbuf_div8_50 : _GEN_8198; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8200 = 6'h33 == _T_498[5:0] ? pgbuf_div8_51 : _GEN_8199; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8201 = 6'h34 == _T_498[5:0] ? pgbuf_div8_52 : _GEN_8200; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8202 = 6'h35 == _T_498[5:0] ? pgbuf_div8_53 : _GEN_8201; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8203 = 6'h36 == _T_498[5:0] ? pgbuf_div8_54 : _GEN_8202; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8204 = 6'h37 == _T_498[5:0] ? pgbuf_div8_55 : _GEN_8203; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8205 = 6'h38 == _T_498[5:0] ? pgbuf_div8_56 : _GEN_8204; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8206 = 6'h39 == _T_498[5:0] ? pgbuf_div8_57 : _GEN_8205; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8207 = 6'h3a == _T_498[5:0] ? pgbuf_div8_58 : _GEN_8206; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8208 = 6'h3b == _T_498[5:0] ? pgbuf_div8_59 : _GEN_8207; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8209 = 6'h3c == _T_498[5:0] ? pgbuf_div8_60 : _GEN_8208; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8210 = 6'h3d == _T_498[5:0] ? pgbuf_div8_61 : _GEN_8209; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8211 = 6'h3e == _T_498[5:0] ? pgbuf_div8_62 : _GEN_8210; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8212 = 6'h3f == _T_498[5:0] ? pgbuf_div8_63 : _GEN_8211; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8145 = 2'h0 == opidx ? _GEN_8212 : _GEN_8132; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8146 = 2'h1 == opidx ? _GEN_8212 : _GEN_8133; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8147 = 2'h2 == opidx ? _GEN_8212 : _GEN_8134; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8148 = 2'h3 == opidx ? _GEN_8212 : _GEN_8135; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8213 = ~_GEN_1128 ? _cnt_T : _GEN_8136; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8214 = cnt[14] ? _GEN_8137 : _GEN_8124; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8215 = cnt[14] ? _GEN_8138 : _GEN_8125; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8216 = cnt[14] ? _GEN_8139 : _GEN_8126; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8217 = cnt[14] ? _GEN_8140 : _GEN_8127; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8218 = cnt[14] ? _GEN_8141 : _GEN_8128; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8219 = cnt[14] ? _GEN_8142 : _GEN_8129; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8220 = cnt[14] ? _GEN_8143 : _GEN_8130; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8221 = cnt[14] ? _GEN_8144 : _GEN_8131; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8222 = cnt[14] ? _GEN_8145 : _GEN_8132; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8223 = cnt[14] ? _GEN_8146 : _GEN_8133; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8224 = cnt[14] ? _GEN_8147 : _GEN_8134; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8225 = cnt[14] ? _GEN_8148 : _GEN_8135; // @[NulCtrlMP.scala 902:29]
  wire [128:0] _GEN_8226 = cnt[14] ? _GEN_8213 : _GEN_8136; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8227 = _GEN_145 | _GEN_8214; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8228 = _GEN_146 | _GEN_8215; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8229 = _GEN_147 | _GEN_8216; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8230 = _GEN_148 | _GEN_8217; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8231 = 2'h0 == opidx ? 5'ha : _GEN_8218; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8232 = 2'h1 == opidx ? 5'ha : _GEN_8219; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8233 = 2'h2 == opidx ? 5'ha : _GEN_8220; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8234 = 2'h3 == opidx ? 5'ha : _GEN_8221; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8240 = 6'h1 == _T_504[5:0] ? pgbuf_div8_1 : pgbuf_div8_0; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8241 = 6'h2 == _T_504[5:0] ? pgbuf_div8_2 : _GEN_8240; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8242 = 6'h3 == _T_504[5:0] ? pgbuf_div8_3 : _GEN_8241; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8243 = 6'h4 == _T_504[5:0] ? pgbuf_div8_4 : _GEN_8242; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8244 = 6'h5 == _T_504[5:0] ? pgbuf_div8_5 : _GEN_8243; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8245 = 6'h6 == _T_504[5:0] ? pgbuf_div8_6 : _GEN_8244; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8246 = 6'h7 == _T_504[5:0] ? pgbuf_div8_7 : _GEN_8245; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8247 = 6'h8 == _T_504[5:0] ? pgbuf_div8_8 : _GEN_8246; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8248 = 6'h9 == _T_504[5:0] ? pgbuf_div8_9 : _GEN_8247; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8249 = 6'ha == _T_504[5:0] ? pgbuf_div8_10 : _GEN_8248; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8250 = 6'hb == _T_504[5:0] ? pgbuf_div8_11 : _GEN_8249; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8251 = 6'hc == _T_504[5:0] ? pgbuf_div8_12 : _GEN_8250; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8252 = 6'hd == _T_504[5:0] ? pgbuf_div8_13 : _GEN_8251; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8253 = 6'he == _T_504[5:0] ? pgbuf_div8_14 : _GEN_8252; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8254 = 6'hf == _T_504[5:0] ? pgbuf_div8_15 : _GEN_8253; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8255 = 6'h10 == _T_504[5:0] ? pgbuf_div8_16 : _GEN_8254; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8256 = 6'h11 == _T_504[5:0] ? pgbuf_div8_17 : _GEN_8255; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8257 = 6'h12 == _T_504[5:0] ? pgbuf_div8_18 : _GEN_8256; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8258 = 6'h13 == _T_504[5:0] ? pgbuf_div8_19 : _GEN_8257; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8259 = 6'h14 == _T_504[5:0] ? pgbuf_div8_20 : _GEN_8258; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8260 = 6'h15 == _T_504[5:0] ? pgbuf_div8_21 : _GEN_8259; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8261 = 6'h16 == _T_504[5:0] ? pgbuf_div8_22 : _GEN_8260; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8262 = 6'h17 == _T_504[5:0] ? pgbuf_div8_23 : _GEN_8261; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8263 = 6'h18 == _T_504[5:0] ? pgbuf_div8_24 : _GEN_8262; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8264 = 6'h19 == _T_504[5:0] ? pgbuf_div8_25 : _GEN_8263; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8265 = 6'h1a == _T_504[5:0] ? pgbuf_div8_26 : _GEN_8264; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8266 = 6'h1b == _T_504[5:0] ? pgbuf_div8_27 : _GEN_8265; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8267 = 6'h1c == _T_504[5:0] ? pgbuf_div8_28 : _GEN_8266; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8268 = 6'h1d == _T_504[5:0] ? pgbuf_div8_29 : _GEN_8267; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8269 = 6'h1e == _T_504[5:0] ? pgbuf_div8_30 : _GEN_8268; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8270 = 6'h1f == _T_504[5:0] ? pgbuf_div8_31 : _GEN_8269; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8271 = 6'h20 == _T_504[5:0] ? pgbuf_div8_32 : _GEN_8270; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8272 = 6'h21 == _T_504[5:0] ? pgbuf_div8_33 : _GEN_8271; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8273 = 6'h22 == _T_504[5:0] ? pgbuf_div8_34 : _GEN_8272; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8274 = 6'h23 == _T_504[5:0] ? pgbuf_div8_35 : _GEN_8273; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8275 = 6'h24 == _T_504[5:0] ? pgbuf_div8_36 : _GEN_8274; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8276 = 6'h25 == _T_504[5:0] ? pgbuf_div8_37 : _GEN_8275; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8277 = 6'h26 == _T_504[5:0] ? pgbuf_div8_38 : _GEN_8276; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8278 = 6'h27 == _T_504[5:0] ? pgbuf_div8_39 : _GEN_8277; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8279 = 6'h28 == _T_504[5:0] ? pgbuf_div8_40 : _GEN_8278; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8280 = 6'h29 == _T_504[5:0] ? pgbuf_div8_41 : _GEN_8279; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8281 = 6'h2a == _T_504[5:0] ? pgbuf_div8_42 : _GEN_8280; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8282 = 6'h2b == _T_504[5:0] ? pgbuf_div8_43 : _GEN_8281; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8283 = 6'h2c == _T_504[5:0] ? pgbuf_div8_44 : _GEN_8282; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8284 = 6'h2d == _T_504[5:0] ? pgbuf_div8_45 : _GEN_8283; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8285 = 6'h2e == _T_504[5:0] ? pgbuf_div8_46 : _GEN_8284; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8286 = 6'h2f == _T_504[5:0] ? pgbuf_div8_47 : _GEN_8285; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8287 = 6'h30 == _T_504[5:0] ? pgbuf_div8_48 : _GEN_8286; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8288 = 6'h31 == _T_504[5:0] ? pgbuf_div8_49 : _GEN_8287; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8289 = 6'h32 == _T_504[5:0] ? pgbuf_div8_50 : _GEN_8288; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8290 = 6'h33 == _T_504[5:0] ? pgbuf_div8_51 : _GEN_8289; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8291 = 6'h34 == _T_504[5:0] ? pgbuf_div8_52 : _GEN_8290; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8292 = 6'h35 == _T_504[5:0] ? pgbuf_div8_53 : _GEN_8291; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8293 = 6'h36 == _T_504[5:0] ? pgbuf_div8_54 : _GEN_8292; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8294 = 6'h37 == _T_504[5:0] ? pgbuf_div8_55 : _GEN_8293; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8295 = 6'h38 == _T_504[5:0] ? pgbuf_div8_56 : _GEN_8294; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8296 = 6'h39 == _T_504[5:0] ? pgbuf_div8_57 : _GEN_8295; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8297 = 6'h3a == _T_504[5:0] ? pgbuf_div8_58 : _GEN_8296; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8298 = 6'h3b == _T_504[5:0] ? pgbuf_div8_59 : _GEN_8297; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8299 = 6'h3c == _T_504[5:0] ? pgbuf_div8_60 : _GEN_8298; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8300 = 6'h3d == _T_504[5:0] ? pgbuf_div8_61 : _GEN_8299; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8301 = 6'h3e == _T_504[5:0] ? pgbuf_div8_62 : _GEN_8300; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8302 = 6'h3f == _T_504[5:0] ? pgbuf_div8_63 : _GEN_8301; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8235 = 2'h0 == opidx ? _GEN_8302 : _GEN_8222; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8236 = 2'h1 == opidx ? _GEN_8302 : _GEN_8223; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8237 = 2'h2 == opidx ? _GEN_8302 : _GEN_8224; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8238 = 2'h3 == opidx ? _GEN_8302 : _GEN_8225; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8303 = ~_GEN_1128 ? _cnt_T : _GEN_8226; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8304 = cnt[15] ? _GEN_8227 : _GEN_8214; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8305 = cnt[15] ? _GEN_8228 : _GEN_8215; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8306 = cnt[15] ? _GEN_8229 : _GEN_8216; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8307 = cnt[15] ? _GEN_8230 : _GEN_8217; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8308 = cnt[15] ? _GEN_8231 : _GEN_8218; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8309 = cnt[15] ? _GEN_8232 : _GEN_8219; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8310 = cnt[15] ? _GEN_8233 : _GEN_8220; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8311 = cnt[15] ? _GEN_8234 : _GEN_8221; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8312 = cnt[15] ? _GEN_8235 : _GEN_8222; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8313 = cnt[15] ? _GEN_8236 : _GEN_8223; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8314 = cnt[15] ? _GEN_8237 : _GEN_8224; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8315 = cnt[15] ? _GEN_8238 : _GEN_8225; // @[NulCtrlMP.scala 902:29]
  wire [128:0] _GEN_8316 = cnt[15] ? _GEN_8303 : _GEN_8226; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8317 = _GEN_145 | _GEN_8304; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8318 = _GEN_146 | _GEN_8305; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8319 = _GEN_147 | _GEN_8306; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8320 = _GEN_148 | _GEN_8307; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8321 = 2'h0 == opidx ? 5'hb : _GEN_8308; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8322 = 2'h1 == opidx ? 5'hb : _GEN_8309; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8323 = 2'h2 == opidx ? 5'hb : _GEN_8310; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8324 = 2'h3 == opidx ? 5'hb : _GEN_8311; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8330 = 6'h1 == _T_510[5:0] ? pgbuf_div8_1 : pgbuf_div8_0; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8331 = 6'h2 == _T_510[5:0] ? pgbuf_div8_2 : _GEN_8330; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8332 = 6'h3 == _T_510[5:0] ? pgbuf_div8_3 : _GEN_8331; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8333 = 6'h4 == _T_510[5:0] ? pgbuf_div8_4 : _GEN_8332; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8334 = 6'h5 == _T_510[5:0] ? pgbuf_div8_5 : _GEN_8333; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8335 = 6'h6 == _T_510[5:0] ? pgbuf_div8_6 : _GEN_8334; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8336 = 6'h7 == _T_510[5:0] ? pgbuf_div8_7 : _GEN_8335; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8337 = 6'h8 == _T_510[5:0] ? pgbuf_div8_8 : _GEN_8336; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8338 = 6'h9 == _T_510[5:0] ? pgbuf_div8_9 : _GEN_8337; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8339 = 6'ha == _T_510[5:0] ? pgbuf_div8_10 : _GEN_8338; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8340 = 6'hb == _T_510[5:0] ? pgbuf_div8_11 : _GEN_8339; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8341 = 6'hc == _T_510[5:0] ? pgbuf_div8_12 : _GEN_8340; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8342 = 6'hd == _T_510[5:0] ? pgbuf_div8_13 : _GEN_8341; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8343 = 6'he == _T_510[5:0] ? pgbuf_div8_14 : _GEN_8342; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8344 = 6'hf == _T_510[5:0] ? pgbuf_div8_15 : _GEN_8343; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8345 = 6'h10 == _T_510[5:0] ? pgbuf_div8_16 : _GEN_8344; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8346 = 6'h11 == _T_510[5:0] ? pgbuf_div8_17 : _GEN_8345; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8347 = 6'h12 == _T_510[5:0] ? pgbuf_div8_18 : _GEN_8346; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8348 = 6'h13 == _T_510[5:0] ? pgbuf_div8_19 : _GEN_8347; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8349 = 6'h14 == _T_510[5:0] ? pgbuf_div8_20 : _GEN_8348; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8350 = 6'h15 == _T_510[5:0] ? pgbuf_div8_21 : _GEN_8349; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8351 = 6'h16 == _T_510[5:0] ? pgbuf_div8_22 : _GEN_8350; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8352 = 6'h17 == _T_510[5:0] ? pgbuf_div8_23 : _GEN_8351; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8353 = 6'h18 == _T_510[5:0] ? pgbuf_div8_24 : _GEN_8352; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8354 = 6'h19 == _T_510[5:0] ? pgbuf_div8_25 : _GEN_8353; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8355 = 6'h1a == _T_510[5:0] ? pgbuf_div8_26 : _GEN_8354; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8356 = 6'h1b == _T_510[5:0] ? pgbuf_div8_27 : _GEN_8355; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8357 = 6'h1c == _T_510[5:0] ? pgbuf_div8_28 : _GEN_8356; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8358 = 6'h1d == _T_510[5:0] ? pgbuf_div8_29 : _GEN_8357; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8359 = 6'h1e == _T_510[5:0] ? pgbuf_div8_30 : _GEN_8358; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8360 = 6'h1f == _T_510[5:0] ? pgbuf_div8_31 : _GEN_8359; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8361 = 6'h20 == _T_510[5:0] ? pgbuf_div8_32 : _GEN_8360; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8362 = 6'h21 == _T_510[5:0] ? pgbuf_div8_33 : _GEN_8361; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8363 = 6'h22 == _T_510[5:0] ? pgbuf_div8_34 : _GEN_8362; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8364 = 6'h23 == _T_510[5:0] ? pgbuf_div8_35 : _GEN_8363; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8365 = 6'h24 == _T_510[5:0] ? pgbuf_div8_36 : _GEN_8364; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8366 = 6'h25 == _T_510[5:0] ? pgbuf_div8_37 : _GEN_8365; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8367 = 6'h26 == _T_510[5:0] ? pgbuf_div8_38 : _GEN_8366; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8368 = 6'h27 == _T_510[5:0] ? pgbuf_div8_39 : _GEN_8367; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8369 = 6'h28 == _T_510[5:0] ? pgbuf_div8_40 : _GEN_8368; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8370 = 6'h29 == _T_510[5:0] ? pgbuf_div8_41 : _GEN_8369; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8371 = 6'h2a == _T_510[5:0] ? pgbuf_div8_42 : _GEN_8370; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8372 = 6'h2b == _T_510[5:0] ? pgbuf_div8_43 : _GEN_8371; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8373 = 6'h2c == _T_510[5:0] ? pgbuf_div8_44 : _GEN_8372; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8374 = 6'h2d == _T_510[5:0] ? pgbuf_div8_45 : _GEN_8373; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8375 = 6'h2e == _T_510[5:0] ? pgbuf_div8_46 : _GEN_8374; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8376 = 6'h2f == _T_510[5:0] ? pgbuf_div8_47 : _GEN_8375; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8377 = 6'h30 == _T_510[5:0] ? pgbuf_div8_48 : _GEN_8376; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8378 = 6'h31 == _T_510[5:0] ? pgbuf_div8_49 : _GEN_8377; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8379 = 6'h32 == _T_510[5:0] ? pgbuf_div8_50 : _GEN_8378; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8380 = 6'h33 == _T_510[5:0] ? pgbuf_div8_51 : _GEN_8379; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8381 = 6'h34 == _T_510[5:0] ? pgbuf_div8_52 : _GEN_8380; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8382 = 6'h35 == _T_510[5:0] ? pgbuf_div8_53 : _GEN_8381; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8383 = 6'h36 == _T_510[5:0] ? pgbuf_div8_54 : _GEN_8382; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8384 = 6'h37 == _T_510[5:0] ? pgbuf_div8_55 : _GEN_8383; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8385 = 6'h38 == _T_510[5:0] ? pgbuf_div8_56 : _GEN_8384; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8386 = 6'h39 == _T_510[5:0] ? pgbuf_div8_57 : _GEN_8385; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8387 = 6'h3a == _T_510[5:0] ? pgbuf_div8_58 : _GEN_8386; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8388 = 6'h3b == _T_510[5:0] ? pgbuf_div8_59 : _GEN_8387; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8389 = 6'h3c == _T_510[5:0] ? pgbuf_div8_60 : _GEN_8388; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8390 = 6'h3d == _T_510[5:0] ? pgbuf_div8_61 : _GEN_8389; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8391 = 6'h3e == _T_510[5:0] ? pgbuf_div8_62 : _GEN_8390; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8392 = 6'h3f == _T_510[5:0] ? pgbuf_div8_63 : _GEN_8391; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8325 = 2'h0 == opidx ? _GEN_8392 : _GEN_8312; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8326 = 2'h1 == opidx ? _GEN_8392 : _GEN_8313; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8327 = 2'h2 == opidx ? _GEN_8392 : _GEN_8314; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8328 = 2'h3 == opidx ? _GEN_8392 : _GEN_8315; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8393 = ~_GEN_1128 ? _cnt_T : _GEN_8316; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8394 = cnt[16] ? _GEN_8317 : _GEN_8304; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8395 = cnt[16] ? _GEN_8318 : _GEN_8305; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8396 = cnt[16] ? _GEN_8319 : _GEN_8306; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8397 = cnt[16] ? _GEN_8320 : _GEN_8307; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8398 = cnt[16] ? _GEN_8321 : _GEN_8308; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8399 = cnt[16] ? _GEN_8322 : _GEN_8309; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8400 = cnt[16] ? _GEN_8323 : _GEN_8310; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8401 = cnt[16] ? _GEN_8324 : _GEN_8311; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8402 = cnt[16] ? _GEN_8325 : _GEN_8312; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8403 = cnt[16] ? _GEN_8326 : _GEN_8313; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8404 = cnt[16] ? _GEN_8327 : _GEN_8314; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8405 = cnt[16] ? _GEN_8328 : _GEN_8315; // @[NulCtrlMP.scala 902:29]
  wire [128:0] _GEN_8406 = cnt[16] ? _GEN_8393 : _GEN_8316; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8407 = _GEN_145 | _GEN_8394; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8408 = _GEN_146 | _GEN_8395; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8409 = _GEN_147 | _GEN_8396; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8410 = _GEN_148 | _GEN_8397; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8411 = 2'h0 == opidx ? 5'hc : _GEN_8398; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8412 = 2'h1 == opidx ? 5'hc : _GEN_8399; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8413 = 2'h2 == opidx ? 5'hc : _GEN_8400; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8414 = 2'h3 == opidx ? 5'hc : _GEN_8401; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8420 = 6'h1 == _T_516[5:0] ? pgbuf_div8_1 : pgbuf_div8_0; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8421 = 6'h2 == _T_516[5:0] ? pgbuf_div8_2 : _GEN_8420; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8422 = 6'h3 == _T_516[5:0] ? pgbuf_div8_3 : _GEN_8421; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8423 = 6'h4 == _T_516[5:0] ? pgbuf_div8_4 : _GEN_8422; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8424 = 6'h5 == _T_516[5:0] ? pgbuf_div8_5 : _GEN_8423; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8425 = 6'h6 == _T_516[5:0] ? pgbuf_div8_6 : _GEN_8424; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8426 = 6'h7 == _T_516[5:0] ? pgbuf_div8_7 : _GEN_8425; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8427 = 6'h8 == _T_516[5:0] ? pgbuf_div8_8 : _GEN_8426; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8428 = 6'h9 == _T_516[5:0] ? pgbuf_div8_9 : _GEN_8427; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8429 = 6'ha == _T_516[5:0] ? pgbuf_div8_10 : _GEN_8428; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8430 = 6'hb == _T_516[5:0] ? pgbuf_div8_11 : _GEN_8429; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8431 = 6'hc == _T_516[5:0] ? pgbuf_div8_12 : _GEN_8430; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8432 = 6'hd == _T_516[5:0] ? pgbuf_div8_13 : _GEN_8431; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8433 = 6'he == _T_516[5:0] ? pgbuf_div8_14 : _GEN_8432; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8434 = 6'hf == _T_516[5:0] ? pgbuf_div8_15 : _GEN_8433; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8435 = 6'h10 == _T_516[5:0] ? pgbuf_div8_16 : _GEN_8434; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8436 = 6'h11 == _T_516[5:0] ? pgbuf_div8_17 : _GEN_8435; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8437 = 6'h12 == _T_516[5:0] ? pgbuf_div8_18 : _GEN_8436; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8438 = 6'h13 == _T_516[5:0] ? pgbuf_div8_19 : _GEN_8437; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8439 = 6'h14 == _T_516[5:0] ? pgbuf_div8_20 : _GEN_8438; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8440 = 6'h15 == _T_516[5:0] ? pgbuf_div8_21 : _GEN_8439; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8441 = 6'h16 == _T_516[5:0] ? pgbuf_div8_22 : _GEN_8440; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8442 = 6'h17 == _T_516[5:0] ? pgbuf_div8_23 : _GEN_8441; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8443 = 6'h18 == _T_516[5:0] ? pgbuf_div8_24 : _GEN_8442; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8444 = 6'h19 == _T_516[5:0] ? pgbuf_div8_25 : _GEN_8443; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8445 = 6'h1a == _T_516[5:0] ? pgbuf_div8_26 : _GEN_8444; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8446 = 6'h1b == _T_516[5:0] ? pgbuf_div8_27 : _GEN_8445; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8447 = 6'h1c == _T_516[5:0] ? pgbuf_div8_28 : _GEN_8446; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8448 = 6'h1d == _T_516[5:0] ? pgbuf_div8_29 : _GEN_8447; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8449 = 6'h1e == _T_516[5:0] ? pgbuf_div8_30 : _GEN_8448; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8450 = 6'h1f == _T_516[5:0] ? pgbuf_div8_31 : _GEN_8449; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8451 = 6'h20 == _T_516[5:0] ? pgbuf_div8_32 : _GEN_8450; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8452 = 6'h21 == _T_516[5:0] ? pgbuf_div8_33 : _GEN_8451; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8453 = 6'h22 == _T_516[5:0] ? pgbuf_div8_34 : _GEN_8452; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8454 = 6'h23 == _T_516[5:0] ? pgbuf_div8_35 : _GEN_8453; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8455 = 6'h24 == _T_516[5:0] ? pgbuf_div8_36 : _GEN_8454; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8456 = 6'h25 == _T_516[5:0] ? pgbuf_div8_37 : _GEN_8455; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8457 = 6'h26 == _T_516[5:0] ? pgbuf_div8_38 : _GEN_8456; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8458 = 6'h27 == _T_516[5:0] ? pgbuf_div8_39 : _GEN_8457; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8459 = 6'h28 == _T_516[5:0] ? pgbuf_div8_40 : _GEN_8458; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8460 = 6'h29 == _T_516[5:0] ? pgbuf_div8_41 : _GEN_8459; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8461 = 6'h2a == _T_516[5:0] ? pgbuf_div8_42 : _GEN_8460; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8462 = 6'h2b == _T_516[5:0] ? pgbuf_div8_43 : _GEN_8461; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8463 = 6'h2c == _T_516[5:0] ? pgbuf_div8_44 : _GEN_8462; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8464 = 6'h2d == _T_516[5:0] ? pgbuf_div8_45 : _GEN_8463; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8465 = 6'h2e == _T_516[5:0] ? pgbuf_div8_46 : _GEN_8464; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8466 = 6'h2f == _T_516[5:0] ? pgbuf_div8_47 : _GEN_8465; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8467 = 6'h30 == _T_516[5:0] ? pgbuf_div8_48 : _GEN_8466; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8468 = 6'h31 == _T_516[5:0] ? pgbuf_div8_49 : _GEN_8467; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8469 = 6'h32 == _T_516[5:0] ? pgbuf_div8_50 : _GEN_8468; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8470 = 6'h33 == _T_516[5:0] ? pgbuf_div8_51 : _GEN_8469; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8471 = 6'h34 == _T_516[5:0] ? pgbuf_div8_52 : _GEN_8470; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8472 = 6'h35 == _T_516[5:0] ? pgbuf_div8_53 : _GEN_8471; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8473 = 6'h36 == _T_516[5:0] ? pgbuf_div8_54 : _GEN_8472; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8474 = 6'h37 == _T_516[5:0] ? pgbuf_div8_55 : _GEN_8473; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8475 = 6'h38 == _T_516[5:0] ? pgbuf_div8_56 : _GEN_8474; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8476 = 6'h39 == _T_516[5:0] ? pgbuf_div8_57 : _GEN_8475; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8477 = 6'h3a == _T_516[5:0] ? pgbuf_div8_58 : _GEN_8476; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8478 = 6'h3b == _T_516[5:0] ? pgbuf_div8_59 : _GEN_8477; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8479 = 6'h3c == _T_516[5:0] ? pgbuf_div8_60 : _GEN_8478; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8480 = 6'h3d == _T_516[5:0] ? pgbuf_div8_61 : _GEN_8479; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8481 = 6'h3e == _T_516[5:0] ? pgbuf_div8_62 : _GEN_8480; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8482 = 6'h3f == _T_516[5:0] ? pgbuf_div8_63 : _GEN_8481; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8415 = 2'h0 == opidx ? _GEN_8482 : _GEN_8402; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8416 = 2'h1 == opidx ? _GEN_8482 : _GEN_8403; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8417 = 2'h2 == opidx ? _GEN_8482 : _GEN_8404; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8418 = 2'h3 == opidx ? _GEN_8482 : _GEN_8405; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8483 = ~_GEN_1128 ? _cnt_T : _GEN_8406; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8484 = cnt[17] ? _GEN_8407 : _GEN_8394; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8485 = cnt[17] ? _GEN_8408 : _GEN_8395; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8486 = cnt[17] ? _GEN_8409 : _GEN_8396; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8487 = cnt[17] ? _GEN_8410 : _GEN_8397; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8488 = cnt[17] ? _GEN_8411 : _GEN_8398; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8489 = cnt[17] ? _GEN_8412 : _GEN_8399; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8490 = cnt[17] ? _GEN_8413 : _GEN_8400; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8491 = cnt[17] ? _GEN_8414 : _GEN_8401; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8492 = cnt[17] ? _GEN_8415 : _GEN_8402; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8493 = cnt[17] ? _GEN_8416 : _GEN_8403; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8494 = cnt[17] ? _GEN_8417 : _GEN_8404; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8495 = cnt[17] ? _GEN_8418 : _GEN_8405; // @[NulCtrlMP.scala 902:29]
  wire [128:0] _GEN_8496 = cnt[17] ? _GEN_8483 : _GEN_8406; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8497 = _GEN_145 | _GEN_8484; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8498 = _GEN_146 | _GEN_8485; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8499 = _GEN_147 | _GEN_8486; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8500 = _GEN_148 | _GEN_8487; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8501 = 2'h0 == opidx ? 5'hd : _GEN_8488; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8502 = 2'h1 == opidx ? 5'hd : _GEN_8489; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8503 = 2'h2 == opidx ? 5'hd : _GEN_8490; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8504 = 2'h3 == opidx ? 5'hd : _GEN_8491; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8510 = 6'h1 == _T_522[5:0] ? pgbuf_div8_1 : pgbuf_div8_0; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8511 = 6'h2 == _T_522[5:0] ? pgbuf_div8_2 : _GEN_8510; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8512 = 6'h3 == _T_522[5:0] ? pgbuf_div8_3 : _GEN_8511; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8513 = 6'h4 == _T_522[5:0] ? pgbuf_div8_4 : _GEN_8512; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8514 = 6'h5 == _T_522[5:0] ? pgbuf_div8_5 : _GEN_8513; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8515 = 6'h6 == _T_522[5:0] ? pgbuf_div8_6 : _GEN_8514; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8516 = 6'h7 == _T_522[5:0] ? pgbuf_div8_7 : _GEN_8515; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8517 = 6'h8 == _T_522[5:0] ? pgbuf_div8_8 : _GEN_8516; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8518 = 6'h9 == _T_522[5:0] ? pgbuf_div8_9 : _GEN_8517; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8519 = 6'ha == _T_522[5:0] ? pgbuf_div8_10 : _GEN_8518; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8520 = 6'hb == _T_522[5:0] ? pgbuf_div8_11 : _GEN_8519; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8521 = 6'hc == _T_522[5:0] ? pgbuf_div8_12 : _GEN_8520; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8522 = 6'hd == _T_522[5:0] ? pgbuf_div8_13 : _GEN_8521; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8523 = 6'he == _T_522[5:0] ? pgbuf_div8_14 : _GEN_8522; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8524 = 6'hf == _T_522[5:0] ? pgbuf_div8_15 : _GEN_8523; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8525 = 6'h10 == _T_522[5:0] ? pgbuf_div8_16 : _GEN_8524; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8526 = 6'h11 == _T_522[5:0] ? pgbuf_div8_17 : _GEN_8525; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8527 = 6'h12 == _T_522[5:0] ? pgbuf_div8_18 : _GEN_8526; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8528 = 6'h13 == _T_522[5:0] ? pgbuf_div8_19 : _GEN_8527; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8529 = 6'h14 == _T_522[5:0] ? pgbuf_div8_20 : _GEN_8528; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8530 = 6'h15 == _T_522[5:0] ? pgbuf_div8_21 : _GEN_8529; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8531 = 6'h16 == _T_522[5:0] ? pgbuf_div8_22 : _GEN_8530; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8532 = 6'h17 == _T_522[5:0] ? pgbuf_div8_23 : _GEN_8531; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8533 = 6'h18 == _T_522[5:0] ? pgbuf_div8_24 : _GEN_8532; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8534 = 6'h19 == _T_522[5:0] ? pgbuf_div8_25 : _GEN_8533; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8535 = 6'h1a == _T_522[5:0] ? pgbuf_div8_26 : _GEN_8534; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8536 = 6'h1b == _T_522[5:0] ? pgbuf_div8_27 : _GEN_8535; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8537 = 6'h1c == _T_522[5:0] ? pgbuf_div8_28 : _GEN_8536; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8538 = 6'h1d == _T_522[5:0] ? pgbuf_div8_29 : _GEN_8537; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8539 = 6'h1e == _T_522[5:0] ? pgbuf_div8_30 : _GEN_8538; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8540 = 6'h1f == _T_522[5:0] ? pgbuf_div8_31 : _GEN_8539; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8541 = 6'h20 == _T_522[5:0] ? pgbuf_div8_32 : _GEN_8540; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8542 = 6'h21 == _T_522[5:0] ? pgbuf_div8_33 : _GEN_8541; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8543 = 6'h22 == _T_522[5:0] ? pgbuf_div8_34 : _GEN_8542; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8544 = 6'h23 == _T_522[5:0] ? pgbuf_div8_35 : _GEN_8543; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8545 = 6'h24 == _T_522[5:0] ? pgbuf_div8_36 : _GEN_8544; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8546 = 6'h25 == _T_522[5:0] ? pgbuf_div8_37 : _GEN_8545; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8547 = 6'h26 == _T_522[5:0] ? pgbuf_div8_38 : _GEN_8546; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8548 = 6'h27 == _T_522[5:0] ? pgbuf_div8_39 : _GEN_8547; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8549 = 6'h28 == _T_522[5:0] ? pgbuf_div8_40 : _GEN_8548; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8550 = 6'h29 == _T_522[5:0] ? pgbuf_div8_41 : _GEN_8549; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8551 = 6'h2a == _T_522[5:0] ? pgbuf_div8_42 : _GEN_8550; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8552 = 6'h2b == _T_522[5:0] ? pgbuf_div8_43 : _GEN_8551; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8553 = 6'h2c == _T_522[5:0] ? pgbuf_div8_44 : _GEN_8552; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8554 = 6'h2d == _T_522[5:0] ? pgbuf_div8_45 : _GEN_8553; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8555 = 6'h2e == _T_522[5:0] ? pgbuf_div8_46 : _GEN_8554; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8556 = 6'h2f == _T_522[5:0] ? pgbuf_div8_47 : _GEN_8555; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8557 = 6'h30 == _T_522[5:0] ? pgbuf_div8_48 : _GEN_8556; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8558 = 6'h31 == _T_522[5:0] ? pgbuf_div8_49 : _GEN_8557; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8559 = 6'h32 == _T_522[5:0] ? pgbuf_div8_50 : _GEN_8558; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8560 = 6'h33 == _T_522[5:0] ? pgbuf_div8_51 : _GEN_8559; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8561 = 6'h34 == _T_522[5:0] ? pgbuf_div8_52 : _GEN_8560; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8562 = 6'h35 == _T_522[5:0] ? pgbuf_div8_53 : _GEN_8561; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8563 = 6'h36 == _T_522[5:0] ? pgbuf_div8_54 : _GEN_8562; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8564 = 6'h37 == _T_522[5:0] ? pgbuf_div8_55 : _GEN_8563; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8565 = 6'h38 == _T_522[5:0] ? pgbuf_div8_56 : _GEN_8564; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8566 = 6'h39 == _T_522[5:0] ? pgbuf_div8_57 : _GEN_8565; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8567 = 6'h3a == _T_522[5:0] ? pgbuf_div8_58 : _GEN_8566; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8568 = 6'h3b == _T_522[5:0] ? pgbuf_div8_59 : _GEN_8567; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8569 = 6'h3c == _T_522[5:0] ? pgbuf_div8_60 : _GEN_8568; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8570 = 6'h3d == _T_522[5:0] ? pgbuf_div8_61 : _GEN_8569; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8571 = 6'h3e == _T_522[5:0] ? pgbuf_div8_62 : _GEN_8570; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8572 = 6'h3f == _T_522[5:0] ? pgbuf_div8_63 : _GEN_8571; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8505 = 2'h0 == opidx ? _GEN_8572 : _GEN_8492; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8506 = 2'h1 == opidx ? _GEN_8572 : _GEN_8493; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8507 = 2'h2 == opidx ? _GEN_8572 : _GEN_8494; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8508 = 2'h3 == opidx ? _GEN_8572 : _GEN_8495; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8573 = ~_GEN_1128 ? _cnt_T : _GEN_8496; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8574 = cnt[18] ? _GEN_8497 : _GEN_8484; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8575 = cnt[18] ? _GEN_8498 : _GEN_8485; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8576 = cnt[18] ? _GEN_8499 : _GEN_8486; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8577 = cnt[18] ? _GEN_8500 : _GEN_8487; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8578 = cnt[18] ? _GEN_8501 : _GEN_8488; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8579 = cnt[18] ? _GEN_8502 : _GEN_8489; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8580 = cnt[18] ? _GEN_8503 : _GEN_8490; // @[NulCtrlMP.scala 902:29]
  wire [4:0] _GEN_8581 = cnt[18] ? _GEN_8504 : _GEN_8491; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8582 = cnt[18] ? _GEN_8505 : _GEN_8492; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8583 = cnt[18] ? _GEN_8506 : _GEN_8493; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8584 = cnt[18] ? _GEN_8507 : _GEN_8494; // @[NulCtrlMP.scala 902:29]
  wire [63:0] _GEN_8585 = cnt[18] ? _GEN_8508 : _GEN_8495; // @[NulCtrlMP.scala 902:29]
  wire [128:0] _GEN_8586 = cnt[18] ? _GEN_8573 : _GEN_8496; // @[NulCtrlMP.scala 902:29]
  wire  _GEN_8587 = _GEN_145 | _GEN_7367; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8588 = _GEN_146 | _GEN_7368; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8589 = _GEN_147 | _GEN_7369; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8590 = _GEN_148 | _GEN_7370; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8591 = 2'h0 == opidx ? 32'h62b023 : _GEN_7371; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8592 = 2'h1 == opidx ? 32'h62b023 : _GEN_7372; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8593 = 2'h2 == opidx ? 32'h62b023 : _GEN_7373; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8594 = 2'h3 == opidx ? 32'h62b023 : _GEN_7374; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8595 = _GEN_1180 ? _cnt_T : _GEN_8586; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8596 = cnt[19] ? _GEN_8587 : _GEN_7367; // @[NulCtrlMP.scala 904:23]
  wire  _GEN_8597 = cnt[19] ? _GEN_8588 : _GEN_7368; // @[NulCtrlMP.scala 904:23]
  wire  _GEN_8598 = cnt[19] ? _GEN_8589 : _GEN_7369; // @[NulCtrlMP.scala 904:23]
  wire  _GEN_8599 = cnt[19] ? _GEN_8590 : _GEN_7370; // @[NulCtrlMP.scala 904:23]
  wire [31:0] _GEN_8600 = cnt[19] ? _GEN_8591 : _GEN_7371; // @[NulCtrlMP.scala 904:23]
  wire [31:0] _GEN_8601 = cnt[19] ? _GEN_8592 : _GEN_7372; // @[NulCtrlMP.scala 904:23]
  wire [31:0] _GEN_8602 = cnt[19] ? _GEN_8593 : _GEN_7373; // @[NulCtrlMP.scala 904:23]
  wire [31:0] _GEN_8603 = cnt[19] ? _GEN_8594 : _GEN_7374; // @[NulCtrlMP.scala 904:23]
  wire [128:0] _GEN_8604 = cnt[19] ? _GEN_8595 : _GEN_8586; // @[NulCtrlMP.scala 904:23]
  wire  _GEN_8605 = _GEN_145 | _GEN_8596; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8606 = _GEN_146 | _GEN_8597; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8607 = _GEN_147 | _GEN_8598; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8608 = _GEN_148 | _GEN_8599; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8609 = 2'h0 == opidx ? 32'h72b423 : _GEN_8600; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8610 = 2'h1 == opidx ? 32'h72b423 : _GEN_8601; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8611 = 2'h2 == opidx ? 32'h72b423 : _GEN_8602; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8612 = 2'h3 == opidx ? 32'h72b423 : _GEN_8603; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8613 = _GEN_1180 ? _cnt_T : _GEN_8604; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8614 = cnt[20] ? _GEN_8605 : _GEN_8596; // @[NulCtrlMP.scala 905:23]
  wire  _GEN_8615 = cnt[20] ? _GEN_8606 : _GEN_8597; // @[NulCtrlMP.scala 905:23]
  wire  _GEN_8616 = cnt[20] ? _GEN_8607 : _GEN_8598; // @[NulCtrlMP.scala 905:23]
  wire  _GEN_8617 = cnt[20] ? _GEN_8608 : _GEN_8599; // @[NulCtrlMP.scala 905:23]
  wire [31:0] _GEN_8618 = cnt[20] ? _GEN_8609 : _GEN_8600; // @[NulCtrlMP.scala 905:23]
  wire [31:0] _GEN_8619 = cnt[20] ? _GEN_8610 : _GEN_8601; // @[NulCtrlMP.scala 905:23]
  wire [31:0] _GEN_8620 = cnt[20] ? _GEN_8611 : _GEN_8602; // @[NulCtrlMP.scala 905:23]
  wire [31:0] _GEN_8621 = cnt[20] ? _GEN_8612 : _GEN_8603; // @[NulCtrlMP.scala 905:23]
  wire [128:0] _GEN_8622 = cnt[20] ? _GEN_8613 : _GEN_8604; // @[NulCtrlMP.scala 905:23]
  wire  _GEN_8623 = _GEN_145 | _GEN_8614; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8624 = _GEN_146 | _GEN_8615; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8625 = _GEN_147 | _GEN_8616; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8626 = _GEN_148 | _GEN_8617; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8627 = 2'h0 == opidx ? 32'h82b823 : _GEN_8618; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8628 = 2'h1 == opidx ? 32'h82b823 : _GEN_8619; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8629 = 2'h2 == opidx ? 32'h82b823 : _GEN_8620; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8630 = 2'h3 == opidx ? 32'h82b823 : _GEN_8621; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8631 = _GEN_1180 ? _cnt_T : _GEN_8622; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8632 = cnt[21] ? _GEN_8623 : _GEN_8614; // @[NulCtrlMP.scala 906:23]
  wire  _GEN_8633 = cnt[21] ? _GEN_8624 : _GEN_8615; // @[NulCtrlMP.scala 906:23]
  wire  _GEN_8634 = cnt[21] ? _GEN_8625 : _GEN_8616; // @[NulCtrlMP.scala 906:23]
  wire  _GEN_8635 = cnt[21] ? _GEN_8626 : _GEN_8617; // @[NulCtrlMP.scala 906:23]
  wire [31:0] _GEN_8636 = cnt[21] ? _GEN_8627 : _GEN_8618; // @[NulCtrlMP.scala 906:23]
  wire [31:0] _GEN_8637 = cnt[21] ? _GEN_8628 : _GEN_8619; // @[NulCtrlMP.scala 906:23]
  wire [31:0] _GEN_8638 = cnt[21] ? _GEN_8629 : _GEN_8620; // @[NulCtrlMP.scala 906:23]
  wire [31:0] _GEN_8639 = cnt[21] ? _GEN_8630 : _GEN_8621; // @[NulCtrlMP.scala 906:23]
  wire [128:0] _GEN_8640 = cnt[21] ? _GEN_8631 : _GEN_8622; // @[NulCtrlMP.scala 906:23]
  wire  _GEN_8641 = _GEN_145 | _GEN_8632; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8642 = _GEN_146 | _GEN_8633; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8643 = _GEN_147 | _GEN_8634; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8644 = _GEN_148 | _GEN_8635; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8645 = 2'h0 == opidx ? 32'h92bc23 : _GEN_8636; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8646 = 2'h1 == opidx ? 32'h92bc23 : _GEN_8637; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8647 = 2'h2 == opidx ? 32'h92bc23 : _GEN_8638; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8648 = 2'h3 == opidx ? 32'h92bc23 : _GEN_8639; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8649 = _GEN_1180 ? _cnt_T : _GEN_8640; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8650 = cnt[22] ? _GEN_8641 : _GEN_8632; // @[NulCtrlMP.scala 907:23]
  wire  _GEN_8651 = cnt[22] ? _GEN_8642 : _GEN_8633; // @[NulCtrlMP.scala 907:23]
  wire  _GEN_8652 = cnt[22] ? _GEN_8643 : _GEN_8634; // @[NulCtrlMP.scala 907:23]
  wire  _GEN_8653 = cnt[22] ? _GEN_8644 : _GEN_8635; // @[NulCtrlMP.scala 907:23]
  wire [31:0] _GEN_8654 = cnt[22] ? _GEN_8645 : _GEN_8636; // @[NulCtrlMP.scala 907:23]
  wire [31:0] _GEN_8655 = cnt[22] ? _GEN_8646 : _GEN_8637; // @[NulCtrlMP.scala 907:23]
  wire [31:0] _GEN_8656 = cnt[22] ? _GEN_8647 : _GEN_8638; // @[NulCtrlMP.scala 907:23]
  wire [31:0] _GEN_8657 = cnt[22] ? _GEN_8648 : _GEN_8639; // @[NulCtrlMP.scala 907:23]
  wire [128:0] _GEN_8658 = cnt[22] ? _GEN_8649 : _GEN_8640; // @[NulCtrlMP.scala 907:23]
  wire  _GEN_8659 = _GEN_145 | _GEN_8650; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8660 = _GEN_146 | _GEN_8651; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8661 = _GEN_147 | _GEN_8652; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8662 = _GEN_148 | _GEN_8653; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8663 = 2'h0 == opidx ? 32'h2a2b023 : _GEN_8654; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8664 = 2'h1 == opidx ? 32'h2a2b023 : _GEN_8655; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8665 = 2'h2 == opidx ? 32'h2a2b023 : _GEN_8656; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8666 = 2'h3 == opidx ? 32'h2a2b023 : _GEN_8657; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8667 = _GEN_1180 ? _cnt_T : _GEN_8658; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8668 = cnt[23] ? _GEN_8659 : _GEN_8650; // @[NulCtrlMP.scala 908:23]
  wire  _GEN_8669 = cnt[23] ? _GEN_8660 : _GEN_8651; // @[NulCtrlMP.scala 908:23]
  wire  _GEN_8670 = cnt[23] ? _GEN_8661 : _GEN_8652; // @[NulCtrlMP.scala 908:23]
  wire  _GEN_8671 = cnt[23] ? _GEN_8662 : _GEN_8653; // @[NulCtrlMP.scala 908:23]
  wire [31:0] _GEN_8672 = cnt[23] ? _GEN_8663 : _GEN_8654; // @[NulCtrlMP.scala 908:23]
  wire [31:0] _GEN_8673 = cnt[23] ? _GEN_8664 : _GEN_8655; // @[NulCtrlMP.scala 908:23]
  wire [31:0] _GEN_8674 = cnt[23] ? _GEN_8665 : _GEN_8656; // @[NulCtrlMP.scala 908:23]
  wire [31:0] _GEN_8675 = cnt[23] ? _GEN_8666 : _GEN_8657; // @[NulCtrlMP.scala 908:23]
  wire [128:0] _GEN_8676 = cnt[23] ? _GEN_8667 : _GEN_8658; // @[NulCtrlMP.scala 908:23]
  wire  _GEN_8677 = _GEN_145 | _GEN_8668; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8678 = _GEN_146 | _GEN_8669; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8679 = _GEN_147 | _GEN_8670; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8680 = _GEN_148 | _GEN_8671; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8681 = 2'h0 == opidx ? 32'h2b2b423 : _GEN_8672; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8682 = 2'h1 == opidx ? 32'h2b2b423 : _GEN_8673; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8683 = 2'h2 == opidx ? 32'h2b2b423 : _GEN_8674; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8684 = 2'h3 == opidx ? 32'h2b2b423 : _GEN_8675; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8685 = _GEN_1180 ? _cnt_T : _GEN_8676; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8686 = cnt[24] ? _GEN_8677 : _GEN_8668; // @[NulCtrlMP.scala 909:23]
  wire  _GEN_8687 = cnt[24] ? _GEN_8678 : _GEN_8669; // @[NulCtrlMP.scala 909:23]
  wire  _GEN_8688 = cnt[24] ? _GEN_8679 : _GEN_8670; // @[NulCtrlMP.scala 909:23]
  wire  _GEN_8689 = cnt[24] ? _GEN_8680 : _GEN_8671; // @[NulCtrlMP.scala 909:23]
  wire [31:0] _GEN_8690 = cnt[24] ? _GEN_8681 : _GEN_8672; // @[NulCtrlMP.scala 909:23]
  wire [31:0] _GEN_8691 = cnt[24] ? _GEN_8682 : _GEN_8673; // @[NulCtrlMP.scala 909:23]
  wire [31:0] _GEN_8692 = cnt[24] ? _GEN_8683 : _GEN_8674; // @[NulCtrlMP.scala 909:23]
  wire [31:0] _GEN_8693 = cnt[24] ? _GEN_8684 : _GEN_8675; // @[NulCtrlMP.scala 909:23]
  wire [128:0] _GEN_8694 = cnt[24] ? _GEN_8685 : _GEN_8676; // @[NulCtrlMP.scala 909:23]
  wire  _GEN_8695 = _GEN_145 | _GEN_8686; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8696 = _GEN_146 | _GEN_8687; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8697 = _GEN_147 | _GEN_8688; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8698 = _GEN_148 | _GEN_8689; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8699 = 2'h0 == opidx ? 32'h2c2b823 : _GEN_8690; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8700 = 2'h1 == opidx ? 32'h2c2b823 : _GEN_8691; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8701 = 2'h2 == opidx ? 32'h2c2b823 : _GEN_8692; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8702 = 2'h3 == opidx ? 32'h2c2b823 : _GEN_8693; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8703 = _GEN_1180 ? _cnt_T : _GEN_8694; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8704 = cnt[25] ? _GEN_8695 : _GEN_8686; // @[NulCtrlMP.scala 910:23]
  wire  _GEN_8705 = cnt[25] ? _GEN_8696 : _GEN_8687; // @[NulCtrlMP.scala 910:23]
  wire  _GEN_8706 = cnt[25] ? _GEN_8697 : _GEN_8688; // @[NulCtrlMP.scala 910:23]
  wire  _GEN_8707 = cnt[25] ? _GEN_8698 : _GEN_8689; // @[NulCtrlMP.scala 910:23]
  wire [31:0] _GEN_8708 = cnt[25] ? _GEN_8699 : _GEN_8690; // @[NulCtrlMP.scala 910:23]
  wire [31:0] _GEN_8709 = cnt[25] ? _GEN_8700 : _GEN_8691; // @[NulCtrlMP.scala 910:23]
  wire [31:0] _GEN_8710 = cnt[25] ? _GEN_8701 : _GEN_8692; // @[NulCtrlMP.scala 910:23]
  wire [31:0] _GEN_8711 = cnt[25] ? _GEN_8702 : _GEN_8693; // @[NulCtrlMP.scala 910:23]
  wire [128:0] _GEN_8712 = cnt[25] ? _GEN_8703 : _GEN_8694; // @[NulCtrlMP.scala 910:23]
  wire  _GEN_8713 = _GEN_145 | _GEN_8704; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8714 = _GEN_146 | _GEN_8705; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8715 = _GEN_147 | _GEN_8706; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8716 = _GEN_148 | _GEN_8707; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8717 = 2'h0 == opidx ? 32'h2d2bc23 : _GEN_8708; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8718 = 2'h1 == opidx ? 32'h2d2bc23 : _GEN_8709; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8719 = 2'h2 == opidx ? 32'h2d2bc23 : _GEN_8710; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8720 = 2'h3 == opidx ? 32'h2d2bc23 : _GEN_8711; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8721 = _GEN_1180 ? _cnt_T : _GEN_8712; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8722 = cnt[26] ? _GEN_8713 : _GEN_8704; // @[NulCtrlMP.scala 911:23]
  wire  _GEN_8723 = cnt[26] ? _GEN_8714 : _GEN_8705; // @[NulCtrlMP.scala 911:23]
  wire  _GEN_8724 = cnt[26] ? _GEN_8715 : _GEN_8706; // @[NulCtrlMP.scala 911:23]
  wire  _GEN_8725 = cnt[26] ? _GEN_8716 : _GEN_8707; // @[NulCtrlMP.scala 911:23]
  wire [31:0] _GEN_8726 = cnt[26] ? _GEN_8717 : _GEN_8708; // @[NulCtrlMP.scala 911:23]
  wire [31:0] _GEN_8727 = cnt[26] ? _GEN_8718 : _GEN_8709; // @[NulCtrlMP.scala 911:23]
  wire [31:0] _GEN_8728 = cnt[26] ? _GEN_8719 : _GEN_8710; // @[NulCtrlMP.scala 911:23]
  wire [31:0] _GEN_8729 = cnt[26] ? _GEN_8720 : _GEN_8711; // @[NulCtrlMP.scala 911:23]
  wire [128:0] _GEN_8730 = cnt[26] ? _GEN_8721 : _GEN_8712; // @[NulCtrlMP.scala 911:23]
  wire  _GEN_8731 = _GEN_145 | _GEN_8722; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8732 = _GEN_146 | _GEN_8723; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8733 = _GEN_147 | _GEN_8724; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8734 = _GEN_148 | _GEN_8725; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8735 = 2'h0 == opidx ? 32'h4028293 : _GEN_8726; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8736 = 2'h1 == opidx ? 32'h4028293 : _GEN_8727; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8737 = 2'h2 == opidx ? 32'h4028293 : _GEN_8728; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8738 = 2'h3 == opidx ? 32'h4028293 : _GEN_8729; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8739 = _GEN_1180 ? _cnt_T : _GEN_8730; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8740 = cnt[27] ? _GEN_8731 : _GEN_8722; // @[NulCtrlMP.scala 912:23]
  wire  _GEN_8741 = cnt[27] ? _GEN_8732 : _GEN_8723; // @[NulCtrlMP.scala 912:23]
  wire  _GEN_8742 = cnt[27] ? _GEN_8733 : _GEN_8724; // @[NulCtrlMP.scala 912:23]
  wire  _GEN_8743 = cnt[27] ? _GEN_8734 : _GEN_8725; // @[NulCtrlMP.scala 912:23]
  wire [31:0] _GEN_8744 = cnt[27] ? _GEN_8735 : _GEN_8726; // @[NulCtrlMP.scala 912:23]
  wire [31:0] _GEN_8745 = cnt[27] ? _GEN_8736 : _GEN_8727; // @[NulCtrlMP.scala 912:23]
  wire [31:0] _GEN_8746 = cnt[27] ? _GEN_8737 : _GEN_8728; // @[NulCtrlMP.scala 912:23]
  wire [31:0] _GEN_8747 = cnt[27] ? _GEN_8738 : _GEN_8729; // @[NulCtrlMP.scala 912:23]
  wire [128:0] _GEN_8748 = cnt[27] ? _GEN_8739 : _GEN_8730; // @[NulCtrlMP.scala 912:23]
  wire  _GEN_8749 = _GEN_145 | _GEN_7375; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_8750 = _GEN_146 | _GEN_7376; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_8751 = _GEN_147 | _GEN_7377; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_8752 = _GEN_148 | _GEN_7378; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_8753 = ~_GEN_1252 ? _cnt_T : _GEN_8748; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_8754 = cnt[28] ? _GEN_8749 : _GEN_7375; // @[NulCtrlMP.scala 913:23]
  wire  _GEN_8755 = cnt[28] ? _GEN_8750 : _GEN_7376; // @[NulCtrlMP.scala 913:23]
  wire  _GEN_8756 = cnt[28] ? _GEN_8751 : _GEN_7377; // @[NulCtrlMP.scala 913:23]
  wire  _GEN_8757 = cnt[28] ? _GEN_8752 : _GEN_7378; // @[NulCtrlMP.scala 913:23]
  wire [128:0] _GEN_8758 = cnt[28] ? _GEN_8753 : _GEN_8748; // @[NulCtrlMP.scala 913:23]
  wire [128:0] _GEN_8759 = _T_526 ? _cnt_T : 129'h400; // @[NulCtrlMP.scala 915:43 916:21 918:21]
  wire [128:0] _GEN_8760 = cnt[29] ? _GEN_8759 : _GEN_8758; // @[NulCtrlMP.scala 914:23]
  wire  _GEN_8762 = _GEN_145 | _GEN_8740; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8763 = _GEN_146 | _GEN_8741; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8764 = _GEN_147 | _GEN_8742; // @[NulCtrlMP.scala 394:{24,24}]
  wire  _GEN_8765 = _GEN_148 | _GEN_8743; // @[NulCtrlMP.scala 394:{24,24}]
  wire [31:0] _GEN_8766 = 2'h0 == opidx ? 32'h330000f : _GEN_8744; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8767 = 2'h1 == opidx ? 32'h330000f : _GEN_8745; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8768 = 2'h2 == opidx ? 32'h330000f : _GEN_8746; // @[NulCtrlMP.scala 395:{28,28}]
  wire [31:0] _GEN_8769 = 2'h3 == opidx ? 32'h330000f : _GEN_8747; // @[NulCtrlMP.scala 395:{28,28}]
  wire [128:0] _GEN_8770 = _GEN_1180 ? _cnt_T : _GEN_8760; // @[NulCtrlMP.scala 396:36 397:17]
  wire  _GEN_8771 = cnt[30] ? _GEN_8762 : _GEN_8740; // @[NulCtrlMP.scala 922:23]
  wire  _GEN_8772 = cnt[30] ? _GEN_8763 : _GEN_8741; // @[NulCtrlMP.scala 922:23]
  wire  _GEN_8773 = cnt[30] ? _GEN_8764 : _GEN_8742; // @[NulCtrlMP.scala 922:23]
  wire  _GEN_8774 = cnt[30] ? _GEN_8765 : _GEN_8743; // @[NulCtrlMP.scala 922:23]
  wire [31:0] _GEN_8775 = cnt[30] ? _GEN_8766 : _GEN_8744; // @[NulCtrlMP.scala 922:23]
  wire [31:0] _GEN_8776 = cnt[30] ? _GEN_8767 : _GEN_8745; // @[NulCtrlMP.scala 922:23]
  wire [31:0] _GEN_8777 = cnt[30] ? _GEN_8768 : _GEN_8746; // @[NulCtrlMP.scala 922:23]
  wire [31:0] _GEN_8778 = cnt[30] ? _GEN_8769 : _GEN_8747; // @[NulCtrlMP.scala 922:23]
  wire [128:0] _GEN_8779 = cnt[30] ? _GEN_8770 : _GEN_8760; // @[NulCtrlMP.scala 922:23]
  wire  _GEN_8780 = _GEN_145 | _GEN_8754; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_8781 = _GEN_146 | _GEN_8755; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_8782 = _GEN_147 | _GEN_8756; // @[NulCtrlMP.scala 401:{30,30}]
  wire  _GEN_8783 = _GEN_148 | _GEN_8757; // @[NulCtrlMP.scala 401:{30,30}]
  wire [128:0] _GEN_8784 = ~_GEN_1252 ? _cnt_T : _GEN_8779; // @[NulCtrlMP.scala 402:36 403:17]
  wire  _GEN_8785 = cnt[31] ? _GEN_8780 : _GEN_8754; // @[NulCtrlMP.scala 923:23]
  wire  _GEN_8786 = cnt[31] ? _GEN_8781 : _GEN_8755; // @[NulCtrlMP.scala 923:23]
  wire  _GEN_8787 = cnt[31] ? _GEN_8782 : _GEN_8756; // @[NulCtrlMP.scala 923:23]
  wire  _GEN_8788 = cnt[31] ? _GEN_8783 : _GEN_8757; // @[NulCtrlMP.scala 923:23]
  wire [128:0] _GEN_8789 = cnt[31] ? _GEN_8784 : _GEN_8779; // @[NulCtrlMP.scala 923:23]
  wire  _GEN_8790 = _GEN_145 | _GEN_8574; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8791 = _GEN_146 | _GEN_8575; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8792 = _GEN_147 | _GEN_8576; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8793 = _GEN_148 | _GEN_8577; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8794 = 2'h0 == opidx ? 5'h5 : _GEN_8578; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8795 = 2'h1 == opidx ? 5'h5 : _GEN_8579; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8796 = 2'h2 == opidx ? 5'h5 : _GEN_8580; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8797 = 2'h3 == opidx ? 5'h5 : _GEN_8581; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8798 = 2'h0 == opidx ? regback_0 : _GEN_8582; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8799 = 2'h1 == opidx ? regback_0 : _GEN_8583; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8800 = 2'h2 == opidx ? regback_0 : _GEN_8584; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8801 = 2'h3 == opidx ? regback_0 : _GEN_8585; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8802 = ~_GEN_1128 ? _cnt_T : _GEN_8789; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8803 = cnt[32] ? _GEN_8790 : _GEN_8574; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8804 = cnt[32] ? _GEN_8791 : _GEN_8575; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8805 = cnt[32] ? _GEN_8792 : _GEN_8576; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8806 = cnt[32] ? _GEN_8793 : _GEN_8577; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8807 = cnt[32] ? _GEN_8794 : _GEN_8578; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8808 = cnt[32] ? _GEN_8795 : _GEN_8579; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8809 = cnt[32] ? _GEN_8796 : _GEN_8580; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8810 = cnt[32] ? _GEN_8797 : _GEN_8581; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8811 = cnt[32] ? _GEN_8798 : _GEN_8582; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8812 = cnt[32] ? _GEN_8799 : _GEN_8583; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8813 = cnt[32] ? _GEN_8800 : _GEN_8584; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8814 = cnt[32] ? _GEN_8801 : _GEN_8585; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_8815 = cnt[32] ? _GEN_8802 : _GEN_8789; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8816 = _GEN_145 | _GEN_8803; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8817 = _GEN_146 | _GEN_8804; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8818 = _GEN_147 | _GEN_8805; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8819 = _GEN_148 | _GEN_8806; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8820 = 2'h0 == opidx ? 5'h6 : _GEN_8807; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8821 = 2'h1 == opidx ? 5'h6 : _GEN_8808; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8822 = 2'h2 == opidx ? 5'h6 : _GEN_8809; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8823 = 2'h3 == opidx ? 5'h6 : _GEN_8810; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8824 = 2'h0 == opidx ? regback_1 : _GEN_8811; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8825 = 2'h1 == opidx ? regback_1 : _GEN_8812; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8826 = 2'h2 == opidx ? regback_1 : _GEN_8813; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8827 = 2'h3 == opidx ? regback_1 : _GEN_8814; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8828 = ~_GEN_1128 ? _cnt_T : _GEN_8815; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8829 = cnt[33] ? _GEN_8816 : _GEN_8803; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8830 = cnt[33] ? _GEN_8817 : _GEN_8804; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8831 = cnt[33] ? _GEN_8818 : _GEN_8805; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8832 = cnt[33] ? _GEN_8819 : _GEN_8806; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8833 = cnt[33] ? _GEN_8820 : _GEN_8807; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8834 = cnt[33] ? _GEN_8821 : _GEN_8808; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8835 = cnt[33] ? _GEN_8822 : _GEN_8809; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8836 = cnt[33] ? _GEN_8823 : _GEN_8810; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8837 = cnt[33] ? _GEN_8824 : _GEN_8811; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8838 = cnt[33] ? _GEN_8825 : _GEN_8812; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8839 = cnt[33] ? _GEN_8826 : _GEN_8813; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8840 = cnt[33] ? _GEN_8827 : _GEN_8814; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_8841 = cnt[33] ? _GEN_8828 : _GEN_8815; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8842 = _GEN_145 | _GEN_8829; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8843 = _GEN_146 | _GEN_8830; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8844 = _GEN_147 | _GEN_8831; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8845 = _GEN_148 | _GEN_8832; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8846 = 2'h0 == opidx ? 5'h7 : _GEN_8833; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8847 = 2'h1 == opidx ? 5'h7 : _GEN_8834; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8848 = 2'h2 == opidx ? 5'h7 : _GEN_8835; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8849 = 2'h3 == opidx ? 5'h7 : _GEN_8836; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8850 = 2'h0 == opidx ? regback_2 : _GEN_8837; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8851 = 2'h1 == opidx ? regback_2 : _GEN_8838; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8852 = 2'h2 == opidx ? regback_2 : _GEN_8839; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8853 = 2'h3 == opidx ? regback_2 : _GEN_8840; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8854 = ~_GEN_1128 ? _cnt_T : _GEN_8841; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8855 = cnt[34] ? _GEN_8842 : _GEN_8829; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8856 = cnt[34] ? _GEN_8843 : _GEN_8830; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8857 = cnt[34] ? _GEN_8844 : _GEN_8831; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8858 = cnt[34] ? _GEN_8845 : _GEN_8832; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8859 = cnt[34] ? _GEN_8846 : _GEN_8833; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8860 = cnt[34] ? _GEN_8847 : _GEN_8834; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8861 = cnt[34] ? _GEN_8848 : _GEN_8835; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8862 = cnt[34] ? _GEN_8849 : _GEN_8836; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8863 = cnt[34] ? _GEN_8850 : _GEN_8837; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8864 = cnt[34] ? _GEN_8851 : _GEN_8838; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8865 = cnt[34] ? _GEN_8852 : _GEN_8839; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8866 = cnt[34] ? _GEN_8853 : _GEN_8840; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_8867 = cnt[34] ? _GEN_8854 : _GEN_8841; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8868 = _GEN_145 | _GEN_8855; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8869 = _GEN_146 | _GEN_8856; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8870 = _GEN_147 | _GEN_8857; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8871 = _GEN_148 | _GEN_8858; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8872 = 2'h0 == opidx ? 5'h8 : _GEN_8859; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8873 = 2'h1 == opidx ? 5'h8 : _GEN_8860; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8874 = 2'h2 == opidx ? 5'h8 : _GEN_8861; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8875 = 2'h3 == opidx ? 5'h8 : _GEN_8862; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8876 = 2'h0 == opidx ? regback_3 : _GEN_8863; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8877 = 2'h1 == opidx ? regback_3 : _GEN_8864; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8878 = 2'h2 == opidx ? regback_3 : _GEN_8865; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8879 = 2'h3 == opidx ? regback_3 : _GEN_8866; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8880 = ~_GEN_1128 ? _cnt_T : _GEN_8867; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8881 = cnt[35] ? _GEN_8868 : _GEN_8855; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8882 = cnt[35] ? _GEN_8869 : _GEN_8856; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8883 = cnt[35] ? _GEN_8870 : _GEN_8857; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8884 = cnt[35] ? _GEN_8871 : _GEN_8858; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8885 = cnt[35] ? _GEN_8872 : _GEN_8859; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8886 = cnt[35] ? _GEN_8873 : _GEN_8860; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8887 = cnt[35] ? _GEN_8874 : _GEN_8861; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8888 = cnt[35] ? _GEN_8875 : _GEN_8862; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8889 = cnt[35] ? _GEN_8876 : _GEN_8863; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8890 = cnt[35] ? _GEN_8877 : _GEN_8864; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8891 = cnt[35] ? _GEN_8878 : _GEN_8865; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8892 = cnt[35] ? _GEN_8879 : _GEN_8866; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_8893 = cnt[35] ? _GEN_8880 : _GEN_8867; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8894 = _GEN_145 | _GEN_8881; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8895 = _GEN_146 | _GEN_8882; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8896 = _GEN_147 | _GEN_8883; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8897 = _GEN_148 | _GEN_8884; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8898 = 2'h0 == opidx ? 5'h9 : _GEN_8885; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8899 = 2'h1 == opidx ? 5'h9 : _GEN_8886; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8900 = 2'h2 == opidx ? 5'h9 : _GEN_8887; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8901 = 2'h3 == opidx ? 5'h9 : _GEN_8888; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8902 = 2'h0 == opidx ? regback_4 : _GEN_8889; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8903 = 2'h1 == opidx ? regback_4 : _GEN_8890; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8904 = 2'h2 == opidx ? regback_4 : _GEN_8891; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8905 = 2'h3 == opidx ? regback_4 : _GEN_8892; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8906 = ~_GEN_1128 ? _cnt_T : _GEN_8893; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8907 = cnt[36] ? _GEN_8894 : _GEN_8881; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8908 = cnt[36] ? _GEN_8895 : _GEN_8882; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8909 = cnt[36] ? _GEN_8896 : _GEN_8883; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8910 = cnt[36] ? _GEN_8897 : _GEN_8884; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8911 = cnt[36] ? _GEN_8898 : _GEN_8885; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8912 = cnt[36] ? _GEN_8899 : _GEN_8886; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8913 = cnt[36] ? _GEN_8900 : _GEN_8887; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8914 = cnt[36] ? _GEN_8901 : _GEN_8888; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8915 = cnt[36] ? _GEN_8902 : _GEN_8889; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8916 = cnt[36] ? _GEN_8903 : _GEN_8890; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8917 = cnt[36] ? _GEN_8904 : _GEN_8891; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8918 = cnt[36] ? _GEN_8905 : _GEN_8892; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_8919 = cnt[36] ? _GEN_8906 : _GEN_8893; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8920 = _GEN_145 | _GEN_8907; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8921 = _GEN_146 | _GEN_8908; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8922 = _GEN_147 | _GEN_8909; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8923 = _GEN_148 | _GEN_8910; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8924 = 2'h0 == opidx ? 5'ha : _GEN_8911; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8925 = 2'h1 == opidx ? 5'ha : _GEN_8912; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8926 = 2'h2 == opidx ? 5'ha : _GEN_8913; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8927 = 2'h3 == opidx ? 5'ha : _GEN_8914; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8928 = 2'h0 == opidx ? regback_5 : _GEN_8915; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8929 = 2'h1 == opidx ? regback_5 : _GEN_8916; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8930 = 2'h2 == opidx ? regback_5 : _GEN_8917; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8931 = 2'h3 == opidx ? regback_5 : _GEN_8918; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8932 = ~_GEN_1128 ? _cnt_T : _GEN_8919; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8933 = cnt[37] ? _GEN_8920 : _GEN_8907; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8934 = cnt[37] ? _GEN_8921 : _GEN_8908; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8935 = cnt[37] ? _GEN_8922 : _GEN_8909; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8936 = cnt[37] ? _GEN_8923 : _GEN_8910; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8937 = cnt[37] ? _GEN_8924 : _GEN_8911; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8938 = cnt[37] ? _GEN_8925 : _GEN_8912; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8939 = cnt[37] ? _GEN_8926 : _GEN_8913; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8940 = cnt[37] ? _GEN_8927 : _GEN_8914; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8941 = cnt[37] ? _GEN_8928 : _GEN_8915; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8942 = cnt[37] ? _GEN_8929 : _GEN_8916; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8943 = cnt[37] ? _GEN_8930 : _GEN_8917; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8944 = cnt[37] ? _GEN_8931 : _GEN_8918; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_8945 = cnt[37] ? _GEN_8932 : _GEN_8919; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8946 = _GEN_145 | _GEN_8933; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8947 = _GEN_146 | _GEN_8934; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8948 = _GEN_147 | _GEN_8935; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8949 = _GEN_148 | _GEN_8936; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8950 = 2'h0 == opidx ? 5'hb : _GEN_8937; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8951 = 2'h1 == opidx ? 5'hb : _GEN_8938; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8952 = 2'h2 == opidx ? 5'hb : _GEN_8939; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8953 = 2'h3 == opidx ? 5'hb : _GEN_8940; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8954 = 2'h0 == opidx ? regback_6 : _GEN_8941; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8955 = 2'h1 == opidx ? regback_6 : _GEN_8942; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8956 = 2'h2 == opidx ? regback_6 : _GEN_8943; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8957 = 2'h3 == opidx ? regback_6 : _GEN_8944; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8958 = ~_GEN_1128 ? _cnt_T : _GEN_8945; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8959 = cnt[38] ? _GEN_8946 : _GEN_8933; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8960 = cnt[38] ? _GEN_8947 : _GEN_8934; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8961 = cnt[38] ? _GEN_8948 : _GEN_8935; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8962 = cnt[38] ? _GEN_8949 : _GEN_8936; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8963 = cnt[38] ? _GEN_8950 : _GEN_8937; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8964 = cnt[38] ? _GEN_8951 : _GEN_8938; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8965 = cnt[38] ? _GEN_8952 : _GEN_8939; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8966 = cnt[38] ? _GEN_8953 : _GEN_8940; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8967 = cnt[38] ? _GEN_8954 : _GEN_8941; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8968 = cnt[38] ? _GEN_8955 : _GEN_8942; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8969 = cnt[38] ? _GEN_8956 : _GEN_8943; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8970 = cnt[38] ? _GEN_8957 : _GEN_8944; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_8971 = cnt[38] ? _GEN_8958 : _GEN_8945; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8972 = _GEN_145 | _GEN_8959; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8973 = _GEN_146 | _GEN_8960; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8974 = _GEN_147 | _GEN_8961; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8975 = _GEN_148 | _GEN_8962; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_8976 = 2'h0 == opidx ? 5'hc : _GEN_8963; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8977 = 2'h1 == opidx ? 5'hc : _GEN_8964; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8978 = 2'h2 == opidx ? 5'hc : _GEN_8965; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_8979 = 2'h3 == opidx ? 5'hc : _GEN_8966; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_8980 = 2'h0 == opidx ? regback_7 : _GEN_8967; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8981 = 2'h1 == opidx ? regback_7 : _GEN_8968; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8982 = 2'h2 == opidx ? regback_7 : _GEN_8969; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_8983 = 2'h3 == opidx ? regback_7 : _GEN_8970; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_8984 = ~_GEN_1128 ? _cnt_T : _GEN_8971; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_8985 = cnt[39] ? _GEN_8972 : _GEN_8959; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8986 = cnt[39] ? _GEN_8973 : _GEN_8960; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8987 = cnt[39] ? _GEN_8974 : _GEN_8961; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8988 = cnt[39] ? _GEN_8975 : _GEN_8962; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8989 = cnt[39] ? _GEN_8976 : _GEN_8963; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8990 = cnt[39] ? _GEN_8977 : _GEN_8964; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8991 = cnt[39] ? _GEN_8978 : _GEN_8965; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_8992 = cnt[39] ? _GEN_8979 : _GEN_8966; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8993 = cnt[39] ? _GEN_8980 : _GEN_8967; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8994 = cnt[39] ? _GEN_8981 : _GEN_8968; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8995 = cnt[39] ? _GEN_8982 : _GEN_8969; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_8996 = cnt[39] ? _GEN_8983 : _GEN_8970; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_8997 = cnt[39] ? _GEN_8984 : _GEN_8971; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_8998 = _GEN_145 | _GEN_8985; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_8999 = _GEN_146 | _GEN_8986; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_9000 = _GEN_147 | _GEN_8987; // @[NulCtrlMP.scala 369:{27,27}]
  wire  _GEN_9001 = _GEN_148 | _GEN_8988; // @[NulCtrlMP.scala 369:{27,27}]
  wire [4:0] _GEN_9002 = 2'h0 == opidx ? 5'hd : _GEN_8989; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_9003 = 2'h1 == opidx ? 5'hd : _GEN_8990; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_9004 = 2'h2 == opidx ? 5'hd : _GEN_8991; // @[NulCtrlMP.scala 370:{28,28}]
  wire [4:0] _GEN_9005 = 2'h3 == opidx ? 5'hd : _GEN_8992; // @[NulCtrlMP.scala 370:{28,28}]
  wire [63:0] _GEN_9006 = 2'h0 == opidx ? regback_8 : _GEN_8993; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_9007 = 2'h1 == opidx ? regback_8 : _GEN_8994; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_9008 = 2'h2 == opidx ? regback_8 : _GEN_8995; // @[NulCtrlMP.scala 371:{30,30}]
  wire [63:0] _GEN_9009 = 2'h3 == opidx ? regback_8 : _GEN_8996; // @[NulCtrlMP.scala 371:{30,30}]
  wire [128:0] _GEN_9010 = ~_GEN_1128 ? _cnt_T : _GEN_8997; // @[NulCtrlMP.scala 372:36 373:17]
  wire  _GEN_9011 = cnt[40] ? _GEN_8998 : _GEN_8985; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_9012 = cnt[40] ? _GEN_8999 : _GEN_8986; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_9013 = cnt[40] ? _GEN_9000 : _GEN_8987; // @[NulCtrlMP.scala 413:32]
  wire  _GEN_9014 = cnt[40] ? _GEN_9001 : _GEN_8988; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_9015 = cnt[40] ? _GEN_9002 : _GEN_8989; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_9016 = cnt[40] ? _GEN_9003 : _GEN_8990; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_9017 = cnt[40] ? _GEN_9004 : _GEN_8991; // @[NulCtrlMP.scala 413:32]
  wire [4:0] _GEN_9018 = cnt[40] ? _GEN_9005 : _GEN_8992; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_9019 = cnt[40] ? _GEN_9006 : _GEN_8993; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_9020 = cnt[40] ? _GEN_9007 : _GEN_8994; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_9021 = cnt[40] ? _GEN_9008 : _GEN_8995; // @[NulCtrlMP.scala 413:32]
  wire [63:0] _GEN_9022 = cnt[40] ? _GEN_9009 : _GEN_8996; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_9023 = cnt[40] ? _GEN_9010 : _GEN_8997; // @[NulCtrlMP.scala 413:32]
  wire [128:0] _GEN_9024 = cnt[41] ? 129'h1 : _GEN_9023; // @[NulCtrlMP.scala 925:23 926:17]
  wire [4:0] _GEN_9025 = cnt[41] ? 5'h5 : _GEN_7444; // @[NulCtrlMP.scala 925:23 927:19]
  wire  _GEN_9029 = state == 5'h14 ? _GEN_7446 : _GEN_125; // @[NulCtrlMP.scala 879:32]
  wire [128:0] _GEN_9112 = state == 5'h14 ? _GEN_9024 : _GEN_7347; // @[NulCtrlMP.scala 879:32]
  wire [4:0] _GEN_9143 = state == 5'h14 ? _GEN_9025 : _GEN_7444; // @[NulCtrlMP.scala 879:32]
  wire  _T_672 = io_tx_ready & io_tx_valid; // @[Decoupled.scala 50:35]
  wire [4:0] _GEN_9144 = io_tx_bits == 8'hff ? 5'h5 : _GEN_9143; // @[NulCtrlMP.scala 946:43 947:17]
  wire  _T_674 = io_rx_ready & io_rx_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_9149 = _T_674 | _GEN_1060; // @[NulCtrlMP.scala 953:23 955:19]
  wire  _GEN_9150 = send_hear | _GEN_7357; // @[NulCtrlMP.scala 939:20 941:19]
  wire [7:0] _GEN_9151 = send_hear ? uart_buffer : _GEN_7358; // @[NulCtrlMP.scala 939:20 942:18]
  wire  _GEN_9155 = send_hear ? _GEN_9029 : 1'h1; // @[NulCtrlMP.scala 939:20 952:19]
  wire [63:0] _GEN_10150 = reset ? 64'h0 : _GEN_2784; // @[NulCtrlMP.scala 164:{35,35}]
  wire [128:0] _GEN_10151 = reset ? 129'h1 : _GEN_9112; // @[NulCtrlMP.scala 345:{22,22}]
  Queue event_queue ( // @[NulCtrlMP.scala 76:29]
    .clock(event_queue_clock),
    .reset(event_queue_reset),
    .io_enq_ready(event_queue_io_enq_ready),
    .io_enq_valid(event_queue_io_enq_valid),
    .io_enq_bits(event_queue_io_enq_bits),
    .io_deq_ready(event_queue_io_deq_ready),
    .io_deq_valid(event_queue_io_deq_valid),
    .io_deq_bits(event_queue_io_deq_bits)
  );
  assign io_cpu_0_ext_itr = state == 5'h4 & _GEN_935; // @[NulCtrlMP.scala 232:33 44:27]
  assign io_cpu_0_stop_fetch = cpu_state_0 == 2'h2 | cpu_state_0 == 2'h1 | _T_6; // @[NulCtrlMP.scala 73:91]
  assign io_cpu_0_regacc_rd = state == 5'h14 ? _GEN_7829 : _GEN_7339; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_0_regacc_wt = state == 5'h14 ? _GEN_9011 : _GEN_7359; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_0_regacc_idx = state == 5'h14 ? _GEN_9015 : _GEN_7343; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_0_regacc_wdata = state == 5'h14 ? _GEN_9019 : _GEN_7363; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_0_inst64 = state == 5'h14 ? _GEN_8771 : _GEN_7367; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_0_inst64_raw = state == 5'h14 ? _GEN_8775 : _GEN_7371; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_0_inst64_nowait = state == 5'hb ? _GEN_3100 : _GEN_2799; // @[NulCtrlMP.scala 653:33]
  assign io_cpu_0_inst64_flush = state == 5'h14 ? _GEN_8785 : _GEN_7375; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_1_ext_itr = state == 5'h4 & _GEN_936; // @[NulCtrlMP.scala 232:33 44:27]
  assign io_cpu_1_stop_fetch = cpu_state_1 == 2'h2 | cpu_state_1 == 2'h1 | _T_11; // @[NulCtrlMP.scala 73:91]
  assign io_cpu_1_regacc_rd = state == 5'h14 ? _GEN_7830 : _GEN_7340; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_1_regacc_wt = state == 5'h14 ? _GEN_9012 : _GEN_7360; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_1_regacc_idx = state == 5'h14 ? _GEN_9016 : _GEN_7344; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_1_regacc_wdata = state == 5'h14 ? _GEN_9020 : _GEN_7364; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_1_inst64 = state == 5'h14 ? _GEN_8772 : _GEN_7368; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_1_inst64_raw = state == 5'h14 ? _GEN_8776 : _GEN_7372; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_1_inst64_nowait = state == 5'hb ? _GEN_3101 : _GEN_2800; // @[NulCtrlMP.scala 653:33]
  assign io_cpu_1_inst64_flush = state == 5'h14 ? _GEN_8786 : _GEN_7376; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_2_ext_itr = state == 5'h4 & _GEN_937; // @[NulCtrlMP.scala 232:33 44:27]
  assign io_cpu_2_stop_fetch = cpu_state_2 == 2'h2 | cpu_state_2 == 2'h1 | _T_16; // @[NulCtrlMP.scala 73:91]
  assign io_cpu_2_regacc_rd = state == 5'h14 ? _GEN_7831 : _GEN_7341; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_2_regacc_wt = state == 5'h14 ? _GEN_9013 : _GEN_7361; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_2_regacc_idx = state == 5'h14 ? _GEN_9017 : _GEN_7345; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_2_regacc_wdata = state == 5'h14 ? _GEN_9021 : _GEN_7365; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_2_inst64 = state == 5'h14 ? _GEN_8773 : _GEN_7369; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_2_inst64_raw = state == 5'h14 ? _GEN_8777 : _GEN_7373; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_2_inst64_nowait = state == 5'hb ? _GEN_3102 : _GEN_2801; // @[NulCtrlMP.scala 653:33]
  assign io_cpu_2_inst64_flush = state == 5'h14 ? _GEN_8787 : _GEN_7377; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_3_ext_itr = state == 5'h4 & _GEN_938; // @[NulCtrlMP.scala 232:33 44:27]
  assign io_cpu_3_stop_fetch = cpu_state_3 == 2'h2 | cpu_state_3 == 2'h1 | _T_21; // @[NulCtrlMP.scala 73:91]
  assign io_cpu_3_regacc_rd = state == 5'h14 ? _GEN_7832 : _GEN_7342; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_3_regacc_wt = state == 5'h14 ? _GEN_9014 : _GEN_7362; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_3_regacc_idx = state == 5'h14 ? _GEN_9018 : _GEN_7346; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_3_regacc_wdata = state == 5'h14 ? _GEN_9022 : _GEN_7366; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_3_inst64 = state == 5'h14 ? _GEN_8774 : _GEN_7370; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_3_inst64_raw = state == 5'h14 ? _GEN_8778 : _GEN_7374; // @[NulCtrlMP.scala 879:32]
  assign io_cpu_3_inst64_nowait = state == 5'hb ? _GEN_3103 : _GEN_2802; // @[NulCtrlMP.scala 653:33]
  assign io_cpu_3_inst64_flush = state == 5'h14 ? _GEN_8788 : _GEN_7378; // @[NulCtrlMP.scala 879:32]
  assign io_tx_valid = state == 5'h19 ? _GEN_9150 : _GEN_7357; // @[NulCtrlMP.scala 938:29]
  assign io_tx_bits = state == 5'h19 ? _GEN_9151 : _GEN_7358; // @[NulCtrlMP.scala 938:29]
  assign io_rx_ready = state == 5'h19 ? _GEN_9155 : _GEN_9029; // @[NulCtrlMP.scala 938:29]
  assign io_dbg_sta = {io_dbg_sta_hi,errno}; // @[Cat.scala 31:58]
  assign io_state = {{3'd0}, state}; // @[NulCtrlMP.scala 959:12]
  assign io_cpu_state = {{6'd0}, cpu_state_0}; // @[NulCtrlMP.scala 960:16]
  assign io_opcode = {opoff,opcode}; // @[Cat.scala 31:58]
  assign io_rx_data = io_rx_bits; // @[NulCtrlMP.scala 962:14]
  assign io_buildTime = 64'h19c22b77194; // @[NulCtrlMP.scala 964:16]
  assign io_uart_buf = uart_buffer; // @[NulCtrlMP.scala 966:15]
  assign event_queue_clock = clock;
  assign event_queue_reset = reset;
  assign event_queue_io_enq_valid = cpu_raised_itr_0 | cpu_raised_itr_1 | cpu_raised_itr_2 | cpu_raised_itr_3; // @[NulCtrlMP.scala 77:42]
  assign event_queue_io_enq_bits = _event_idx_T[0] ? 2'h0 : _event_idx_T_6; // @[Mux.scala 47:70]
  assign event_queue_io_deq_ready = state == 5'h8; // @[NulCtrlMP.scala 334:40]
  always @(posedge clock) begin
    if (reset) begin // @[NulCtrlMP.scala 41:28]
      cpu_state_0 <= 2'h0; // @[NulCtrlMP.scala 41:28]
    end else if (state == 5'hb) begin // @[NulCtrlMP.scala 653:33]
      if (cnt[14]) begin // @[NulCtrlMP.scala 685:23]
        if (_GEN_1180) begin // @[NulCtrlMP.scala 688:40]
          cpu_state_0 <= _GEN_3092;
        end else begin
          cpu_state_0 <= _GEN_2803;
        end
      end else begin
        cpu_state_0 <= _GEN_2803;
      end
    end else begin
      cpu_state_0 <= _GEN_2803;
    end
    if (reset) begin // @[NulCtrlMP.scala 41:28]
      cpu_state_1 <= 2'h0; // @[NulCtrlMP.scala 41:28]
    end else if (state == 5'hb) begin // @[NulCtrlMP.scala 653:33]
      if (cnt[14]) begin // @[NulCtrlMP.scala 685:23]
        if (_GEN_1180) begin // @[NulCtrlMP.scala 688:40]
          cpu_state_1 <= _GEN_3093;
        end else begin
          cpu_state_1 <= _GEN_2804;
        end
      end else begin
        cpu_state_1 <= _GEN_2804;
      end
    end else begin
      cpu_state_1 <= _GEN_2804;
    end
    if (reset) begin // @[NulCtrlMP.scala 41:28]
      cpu_state_2 <= 2'h0; // @[NulCtrlMP.scala 41:28]
    end else if (state == 5'hb) begin // @[NulCtrlMP.scala 653:33]
      if (cnt[14]) begin // @[NulCtrlMP.scala 685:23]
        if (_GEN_1180) begin // @[NulCtrlMP.scala 688:40]
          cpu_state_2 <= _GEN_3094;
        end else begin
          cpu_state_2 <= _GEN_2805;
        end
      end else begin
        cpu_state_2 <= _GEN_2805;
      end
    end else begin
      cpu_state_2 <= _GEN_2805;
    end
    if (reset) begin // @[NulCtrlMP.scala 41:28]
      cpu_state_3 <= 2'h0; // @[NulCtrlMP.scala 41:28]
    end else if (state == 5'hb) begin // @[NulCtrlMP.scala 653:33]
      if (cnt[14]) begin // @[NulCtrlMP.scala 685:23]
        if (_GEN_1180) begin // @[NulCtrlMP.scala 688:40]
          cpu_state_3 <= _GEN_3095;
        end else begin
          cpu_state_3 <= _GEN_2806;
        end
      end else begin
        cpu_state_3 <= _GEN_2806;
      end
    end else begin
      cpu_state_3 <= _GEN_2806;
    end
    if (reset) begin // @[NulCtrlMP.scala 55:29]
      global_clk <= 64'h0; // @[NulCtrlMP.scala 55:29]
    end else begin
      global_clk <= _global_clk_T_1; // @[NulCtrlMP.scala 58:16]
    end
    if (reset) begin // @[NulCtrlMP.scala 56:27]
      user_clk_0 <= 64'h0; // @[NulCtrlMP.scala 56:27]
    end else if (io_cpu_0_priv == 2'h0) begin // @[NulCtrlMP.scala 60:38]
      user_clk_0 <= _user_clk_0_T_1; // @[NulCtrlMP.scala 61:25]
    end
    if (reset) begin // @[NulCtrlMP.scala 56:27]
      user_clk_1 <= 64'h0; // @[NulCtrlMP.scala 56:27]
    end else if (io_cpu_1_priv == 2'h0) begin // @[NulCtrlMP.scala 60:38]
      user_clk_1 <= _user_clk_1_T_1; // @[NulCtrlMP.scala 61:25]
    end
    if (reset) begin // @[NulCtrlMP.scala 56:27]
      user_clk_2 <= 64'h0; // @[NulCtrlMP.scala 56:27]
    end else if (io_cpu_2_priv == 2'h0) begin // @[NulCtrlMP.scala 60:38]
      user_clk_2 <= _user_clk_2_T_1; // @[NulCtrlMP.scala 61:25]
    end
    if (reset) begin // @[NulCtrlMP.scala 56:27]
      user_clk_3 <= 64'h0; // @[NulCtrlMP.scala 56:27]
    end else if (io_cpu_3_priv == 2'h0) begin // @[NulCtrlMP.scala 60:38]
      user_clk_3 <= _user_clk_3_T_1; // @[NulCtrlMP.scala 61:25]
    end
    if (reset) begin // @[NulCtrlMP.scala 65:33]
      cpu_raised_itr_0 <= 1'h0; // @[NulCtrlMP.scala 65:33]
    end else if (has_itr & event_queue_io_enq_ready) begin // @[NulCtrlMP.scala 81:47]
      if (2'h0 == event_idx) begin // @[NulCtrlMP.scala 82:35]
        cpu_raised_itr_0 <= 1'h0; // @[NulCtrlMP.scala 82:35]
      end else begin
        cpu_raised_itr_0 <= _GEN_4;
      end
    end else begin
      cpu_raised_itr_0 <= _GEN_4;
    end
    if (reset) begin // @[NulCtrlMP.scala 65:33]
      cpu_raised_itr_1 <= 1'h0; // @[NulCtrlMP.scala 65:33]
    end else if (has_itr & event_queue_io_enq_ready) begin // @[NulCtrlMP.scala 81:47]
      if (2'h1 == event_idx) begin // @[NulCtrlMP.scala 82:35]
        cpu_raised_itr_1 <= 1'h0; // @[NulCtrlMP.scala 82:35]
      end else begin
        cpu_raised_itr_1 <= _GEN_6;
      end
    end else begin
      cpu_raised_itr_1 <= _GEN_6;
    end
    if (reset) begin // @[NulCtrlMP.scala 65:33]
      cpu_raised_itr_2 <= 1'h0; // @[NulCtrlMP.scala 65:33]
    end else if (has_itr & event_queue_io_enq_ready) begin // @[NulCtrlMP.scala 81:47]
      if (2'h2 == event_idx) begin // @[NulCtrlMP.scala 82:35]
        cpu_raised_itr_2 <= 1'h0; // @[NulCtrlMP.scala 82:35]
      end else begin
        cpu_raised_itr_2 <= _GEN_8;
      end
    end else begin
      cpu_raised_itr_2 <= _GEN_8;
    end
    if (reset) begin // @[NulCtrlMP.scala 65:33]
      cpu_raised_itr_3 <= 1'h0; // @[NulCtrlMP.scala 65:33]
    end else if (has_itr & event_queue_io_enq_ready) begin // @[NulCtrlMP.scala 81:47]
      if (2'h3 == event_idx) begin // @[NulCtrlMP.scala 82:35]
        cpu_raised_itr_3 <= 1'h0; // @[NulCtrlMP.scala 82:35]
      end else begin
        cpu_raised_itr_3 <= _GEN_10;
      end
    end else begin
      cpu_raised_itr_3 <= _GEN_10;
    end
    if (reset) begin // @[NulCtrlMP.scala 66:28]
      last_priv_0 <= 2'h3; // @[NulCtrlMP.scala 66:28]
    end else begin
      last_priv_0 <= io_cpu_0_priv; // @[NulCtrlMP.scala 68:22]
    end
    if (reset) begin // @[NulCtrlMP.scala 66:28]
      last_priv_1 <= 2'h3; // @[NulCtrlMP.scala 66:28]
    end else begin
      last_priv_1 <= io_cpu_1_priv; // @[NulCtrlMP.scala 68:22]
    end
    if (reset) begin // @[NulCtrlMP.scala 66:28]
      last_priv_2 <= 2'h3; // @[NulCtrlMP.scala 66:28]
    end else begin
      last_priv_2 <= io_cpu_2_priv; // @[NulCtrlMP.scala 68:22]
    end
    if (reset) begin // @[NulCtrlMP.scala 66:28]
      last_priv_3 <= 2'h3; // @[NulCtrlMP.scala 66:28]
    end else begin
      last_priv_3 <= io_cpu_3_priv; // @[NulCtrlMP.scala 68:22]
    end
    if (reset) begin // @[NulCtrlMP.scala 140:24]
      state <= 5'h0; // @[NulCtrlMP.scala 140:24]
    end else if (state == 5'h19) begin // @[NulCtrlMP.scala 938:29]
      if (send_hear) begin // @[NulCtrlMP.scala 939:20]
        if (_T_672) begin // @[NulCtrlMP.scala 943:23]
          state <= _GEN_9144;
        end else begin
          state <= _GEN_9143;
        end
      end else begin
        state <= _GEN_9143;
      end
    end else begin
      state <= _GEN_9143;
    end
    if (reset) begin // @[NulCtrlMP.scala 141:30]
      trans_bytes <= 10'h0; // @[NulCtrlMP.scala 141:30]
    end else if (state == 5'h6) begin // @[NulCtrlMP.scala 318:36]
      if (io_tx_ready) begin // @[NulCtrlMP.scala 321:27]
        if (_T_70) begin // @[NulCtrlMP.scala 322:51]
          trans_bytes <= 10'h0; // @[NulCtrlMP.scala 324:29]
        end else begin
          trans_bytes <= _GEN_1078;
        end
      end else begin
        trans_bytes <= _GEN_1078;
      end
    end else begin
      trans_bytes <= _GEN_1078;
    end
    if (reset) begin // @[NulCtrlMP.scala 142:28]
      trans_pos <= 10'h0; // @[NulCtrlMP.scala 142:28]
    end else if (state == 5'h6) begin // @[NulCtrlMP.scala 318:36]
      if (io_tx_ready) begin // @[NulCtrlMP.scala 321:27]
        if (_T_69 == trans_bytes) begin // @[NulCtrlMP.scala 222:51]
          trans_pos <= 10'h0; // @[NulCtrlMP.scala 223:27]
        end else begin
          trans_pos <= _T_69; // @[NulCtrlMP.scala 227:27]
        end
      end else begin
        trans_pos <= _GEN_1077;
      end
    end else begin
      trans_pos <= _GEN_1077;
    end
    if (reset) begin // @[NulCtrlMP.scala 144:24]
      errno <= 6'h0; // @[NulCtrlMP.scala 144:24]
    end else if (state == 5'h2) begin // @[NulCtrlMP.scala 180:37]
      if (io_rx_valid) begin // @[NulCtrlMP.scala 182:27]
        if (!(rxop == 5'h1 | rxop == 5'h2 | rxop == 5'h5 | rxop == 5'h7 | rxop == 5'h11 | rxop == 5'h13)) begin // @[NulCtrlMP.scala 190:155]
          errno <= _GEN_70;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 149:25]
      opcode <= 5'h0; // @[NulCtrlMP.scala 149:25]
    end else if (state == 5'h2) begin // @[NulCtrlMP.scala 180:37]
      if (io_rx_valid) begin // @[NulCtrlMP.scala 182:27]
        opcode <= rxop; // @[NulCtrlMP.scala 185:20]
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 150:24]
      opoff <= 3'h0; // @[NulCtrlMP.scala 150:24]
    end else if (state == 5'h2) begin // @[NulCtrlMP.scala 180:37]
      if (io_rx_valid) begin // @[NulCtrlMP.scala 182:27]
        opoff <= rxoff; // @[NulCtrlMP.scala 186:19]
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_1 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h1) begin // @[NulCtrlMP.scala 421:35]
      if (cnt[8]) begin // @[NulCtrlMP.scala 442:22]
        if (init_cnt == 2'h3) begin // @[NulCtrlMP.scala 444:47]
          oparg_1 <= _GEN_1109;
        end else begin
          oparg_1 <= nextidx; // @[NulCtrlMP.scala 448:26]
        end
      end else begin
        oparg_1 <= _GEN_1109;
      end
    end else begin
      oparg_1 <= _GEN_1109;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_2 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      oparg_2 <= _GEN_128;
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'h2 == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_2 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_2 <= _GEN_128;
      end
    end else begin
      oparg_2 <= _GEN_128;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_3 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      oparg_3 <= _GEN_129;
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'h3 == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_3 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_3 <= _GEN_129;
      end
    end else begin
      oparg_3 <= _GEN_129;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_4 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      oparg_4 <= _GEN_130;
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'h4 == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_4 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_4 <= _GEN_130;
      end
    end else begin
      oparg_4 <= _GEN_130;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_5 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      oparg_5 <= _GEN_131;
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'h5 == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_5 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_5 <= _GEN_131;
      end
    end else begin
      oparg_5 <= _GEN_131;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_6 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      oparg_6 <= _GEN_132;
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'h6 == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_6 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_6 <= _GEN_132;
      end
    end else begin
      oparg_6 <= _GEN_132;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_7 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (5'h0 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_7 <= _GEN_133;
      end else if (5'h1 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_7 <= _GEN_133;
      end else begin
        oparg_7 <= _GEN_851;
      end
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'h7 == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_7 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_7 <= _GEN_133;
      end
    end else begin
      oparg_7 <= _GEN_133;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_8 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (5'h0 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_8 <= _GEN_134;
      end else if (5'h1 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_8 <= _GEN_134;
      end else begin
        oparg_8 <= _GEN_852;
      end
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'h8 == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_8 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_8 <= _GEN_134;
      end
    end else begin
      oparg_8 <= _GEN_134;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_9 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (5'h0 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_9 <= _GEN_135;
      end else if (5'h1 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_9 <= _GEN_135;
      end else begin
        oparg_9 <= _GEN_853;
      end
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'h9 == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_9 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_9 <= _GEN_135;
      end
    end else begin
      oparg_9 <= _GEN_135;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_10 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (5'h0 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_10 <= _GEN_136;
      end else if (5'h1 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_10 <= _GEN_136;
      end else begin
        oparg_10 <= _GEN_854;
      end
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'ha == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_10 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_10 <= _GEN_136;
      end
    end else begin
      oparg_10 <= _GEN_136;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_11 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (5'h0 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_11 <= _GEN_137;
      end else if (5'h1 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_11 <= _GEN_137;
      end else begin
        oparg_11 <= _GEN_855;
      end
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'hb == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_11 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_11 <= _GEN_137;
      end
    end else begin
      oparg_11 <= _GEN_137;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_12 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (5'h0 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_12 <= _GEN_138;
      end else if (5'h1 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_12 <= _GEN_138;
      end else begin
        oparg_12 <= _GEN_856;
      end
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'hc == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_12 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_12 <= _GEN_138;
      end
    end else begin
      oparg_12 <= _GEN_138;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_13 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (5'h0 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_13 <= _GEN_139;
      end else if (5'h1 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_13 <= _GEN_139;
      end else begin
        oparg_13 <= _GEN_857;
      end
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'hd == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_13 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_13 <= _GEN_139;
      end
    end else begin
      oparg_13 <= _GEN_139;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_14 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (5'h0 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_14 <= _GEN_140;
      end else if (5'h1 == opcode) begin // @[NulCtrlMP.scala 236:24]
        oparg_14 <= _GEN_140;
      end else begin
        oparg_14 <= _GEN_858;
      end
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'he == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_14 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_14 <= _GEN_140;
      end
    end else begin
      oparg_14 <= _GEN_140;
    end
    if (reset) begin // @[NulCtrlMP.scala 151:24]
      oparg_15 <= 8'h0; // @[NulCtrlMP.scala 151:24]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      oparg_15 <= _GEN_141;
    end else if (_T_66 & io_rx_valid) begin // @[NulCtrlMP.scala 295:57]
      if (4'hf == trans_pos[3:0]) begin // @[NulCtrlMP.scala 296:26]
        oparg_15 <= io_rx_bits; // @[NulCtrlMP.scala 296:26]
      end else begin
        oparg_15 <= _GEN_141;
      end
    end else begin
      oparg_15 <= _GEN_141;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_0 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h10) begin // @[NulCtrlMP.scala 702:33]
      if (cnt[6]) begin // @[NulCtrlMP.scala 708:22]
        if (_T_122) begin // @[NulCtrlMP.scala 361:36]
          retarg_0 <= _GEN_1349[7:0]; // @[NulCtrlMP.scala 364:33]
        end else begin
          retarg_0 <= _GEN_1795;
        end
      end else begin
        retarg_0 <= _GEN_1795;
      end
    end else begin
      retarg_0 <= _GEN_1795;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_1 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h10) begin // @[NulCtrlMP.scala 702:33]
      if (cnt[6]) begin // @[NulCtrlMP.scala 708:22]
        if (_T_122) begin // @[NulCtrlMP.scala 361:36]
          retarg_1 <= _GEN_1349[15:8]; // @[NulCtrlMP.scala 364:33]
        end else begin
          retarg_1 <= _GEN_2452;
        end
      end else begin
        retarg_1 <= _GEN_2452;
      end
    end else begin
      retarg_1 <= _GEN_2452;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_2 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h10) begin // @[NulCtrlMP.scala 702:33]
      if (cnt[6]) begin // @[NulCtrlMP.scala 708:22]
        if (_T_122) begin // @[NulCtrlMP.scala 361:36]
          retarg_2 <= _GEN_1349[23:16]; // @[NulCtrlMP.scala 364:33]
        end else begin
          retarg_2 <= _GEN_2453;
        end
      end else begin
        retarg_2 <= _GEN_2453;
      end
    end else begin
      retarg_2 <= _GEN_2453;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_3 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h10) begin // @[NulCtrlMP.scala 702:33]
      if (cnt[6]) begin // @[NulCtrlMP.scala 708:22]
        if (_T_122) begin // @[NulCtrlMP.scala 361:36]
          retarg_3 <= _GEN_1349[31:24]; // @[NulCtrlMP.scala 364:33]
        end else begin
          retarg_3 <= _GEN_2454;
        end
      end else begin
        retarg_3 <= _GEN_2454;
      end
    end else begin
      retarg_3 <= _GEN_2454;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_4 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h10) begin // @[NulCtrlMP.scala 702:33]
      if (cnt[6]) begin // @[NulCtrlMP.scala 708:22]
        if (_T_122) begin // @[NulCtrlMP.scala 361:36]
          retarg_4 <= _GEN_1349[39:32]; // @[NulCtrlMP.scala 364:33]
        end else begin
          retarg_4 <= _GEN_2455;
        end
      end else begin
        retarg_4 <= _GEN_2455;
      end
    end else begin
      retarg_4 <= _GEN_2455;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_5 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h10) begin // @[NulCtrlMP.scala 702:33]
      if (cnt[6]) begin // @[NulCtrlMP.scala 708:22]
        if (_T_122) begin // @[NulCtrlMP.scala 361:36]
          retarg_5 <= _GEN_1349[47:40]; // @[NulCtrlMP.scala 364:33]
        end else begin
          retarg_5 <= _GEN_2456;
        end
      end else begin
        retarg_5 <= _GEN_2456;
      end
    end else begin
      retarg_5 <= _GEN_2456;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_6 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h10) begin // @[NulCtrlMP.scala 702:33]
      if (cnt[6]) begin // @[NulCtrlMP.scala 708:22]
        if (_T_122) begin // @[NulCtrlMP.scala 361:36]
          retarg_6 <= _GEN_1349[55:48]; // @[NulCtrlMP.scala 364:33]
        end else begin
          retarg_6 <= _GEN_2457;
        end
      end else begin
        retarg_6 <= _GEN_2457;
      end
    end else begin
      retarg_6 <= _GEN_2457;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_7 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h10) begin // @[NulCtrlMP.scala 702:33]
      if (cnt[6]) begin // @[NulCtrlMP.scala 708:22]
        if (_T_122) begin // @[NulCtrlMP.scala 361:36]
          retarg_7 <= _GEN_1349[63:56]; // @[NulCtrlMP.scala 364:33]
        end else begin
          retarg_7 <= _GEN_2458;
        end
      end else begin
        retarg_7 <= _GEN_2458;
      end
    end else begin
      retarg_7 <= _GEN_2458;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_8 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h9) begin // @[NulCtrlMP.scala 569:32]
      if (cnt[14]) begin // @[NulCtrlMP.scala 580:23]
        if (retarg_1 == 8'h8) begin // @[NulCtrlMP.scala 582:46]
          retarg_8 <= regback_0[7:0]; // @[NulCtrlMP.scala 584:33]
        end else begin
          retarg_8 <= _GEN_2309;
        end
      end else begin
        retarg_8 <= _GEN_2309;
      end
    end else begin
      retarg_8 <= _GEN_1941;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_9 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h9) begin // @[NulCtrlMP.scala 569:32]
      if (cnt[14]) begin // @[NulCtrlMP.scala 580:23]
        if (retarg_1 == 8'h8) begin // @[NulCtrlMP.scala 582:46]
          retarg_9 <= regback_0[15:8]; // @[NulCtrlMP.scala 584:33]
        end else begin
          retarg_9 <= _GEN_2310;
        end
      end else begin
        retarg_9 <= _GEN_2310;
      end
    end else begin
      retarg_9 <= _GEN_1942;
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_10 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h9) begin // @[NulCtrlMP.scala 569:32]
      if (cnt[14]) begin // @[NulCtrlMP.scala 580:23]
        if (retarg_1 == 8'h8) begin // @[NulCtrlMP.scala 582:46]
          retarg_10 <= regback_0[23:16]; // @[NulCtrlMP.scala 584:33]
        end else begin
          retarg_10 <= _GEN_2311;
        end
      end else begin
        retarg_10 <= _GEN_2311;
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_11 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h9) begin // @[NulCtrlMP.scala 569:32]
      if (cnt[14]) begin // @[NulCtrlMP.scala 580:23]
        if (retarg_1 == 8'h8) begin // @[NulCtrlMP.scala 582:46]
          retarg_11 <= regback_0[31:24]; // @[NulCtrlMP.scala 584:33]
        end else begin
          retarg_11 <= _GEN_2312;
        end
      end else begin
        retarg_11 <= _GEN_2312;
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_12 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h9) begin // @[NulCtrlMP.scala 569:32]
      if (cnt[14]) begin // @[NulCtrlMP.scala 580:23]
        if (retarg_1 == 8'h8) begin // @[NulCtrlMP.scala 582:46]
          retarg_12 <= regback_0[39:32]; // @[NulCtrlMP.scala 584:33]
        end else begin
          retarg_12 <= _GEN_2313;
        end
      end else begin
        retarg_12 <= _GEN_2313;
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 152:25]
      retarg_13 <= 8'h0; // @[NulCtrlMP.scala 152:25]
    end else if (state == 5'h9) begin // @[NulCtrlMP.scala 569:32]
      if (cnt[14]) begin // @[NulCtrlMP.scala 580:23]
        if (retarg_1 == 8'h8) begin // @[NulCtrlMP.scala 582:46]
          retarg_13 <= regback_0[47:40]; // @[NulCtrlMP.scala 584:33]
        end else begin
          retarg_13 <= _GEN_2314;
        end
      end else begin
        retarg_13 <= _GEN_2314;
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_0_0 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_0_0 <= _GEN_867;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_0_1 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_0_1 <= _GEN_868;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_0_2 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_0_2 <= _GEN_869;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_0_3 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_0_3 <= _GEN_870;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_1_0 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_1_0 <= _GEN_871;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_1_1 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_1_1 <= _GEN_872;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_1_2 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_1_2 <= _GEN_873;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_1_3 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_1_3 <= _GEN_874;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_2_0 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_2_0 <= _GEN_875;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_2_1 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_2_1 <= _GEN_876;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_2_2 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_2_2 <= _GEN_877;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_2_3 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_2_3 <= _GEN_878;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_3_0 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_3_0 <= _GEN_879;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_3_1 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_3_1 <= _GEN_880;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_3_2 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_3_2 <= _GEN_881;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 162:31]
      hfutex_masks_3_3 <= 48'h0; // @[NulCtrlMP.scala 162:31]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_masks_3_3 <= _GEN_882;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 163:29]
      hfutex_pos_0 <= 2'h0; // @[NulCtrlMP.scala 163:29]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_pos_0 <= _GEN_883;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 163:29]
      hfutex_pos_1 <= 2'h0; // @[NulCtrlMP.scala 163:29]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_pos_1 <= _GEN_884;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 163:29]
      hfutex_pos_2 <= 2'h0; // @[NulCtrlMP.scala 163:29]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_pos_2 <= _GEN_885;
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 163:29]
      hfutex_pos_3 <= 2'h0; // @[NulCtrlMP.scala 163:29]
    end else if (state == 5'h4) begin // @[NulCtrlMP.scala 232:33]
      if (!(5'h0 == opcode)) begin // @[NulCtrlMP.scala 236:24]
        if (!(5'h1 == opcode)) begin // @[NulCtrlMP.scala 236:24]
          hfutex_pos_3 <= _GEN_886;
        end
      end
    end
    hfutex_match_reg <= _GEN_10150[47:0]; // @[NulCtrlMP.scala 164:{35,35}]
    if (reset) begin // @[NulCtrlMP.scala 169:28]
      send_hear <= 1'h0; // @[NulCtrlMP.scala 169:28]
    end else if (state == 5'h19) begin // @[NulCtrlMP.scala 938:29]
      if (send_hear) begin // @[NulCtrlMP.scala 939:20]
        if (_T_672) begin // @[NulCtrlMP.scala 943:23]
          send_hear <= 1'h0; // @[NulCtrlMP.scala 944:19]
        end else begin
          send_hear <= _GEN_1060;
        end
      end else begin
        send_hear <= _GEN_9149;
      end
    end else begin
      send_hear <= _GEN_1060;
    end
    if (reset) begin // @[NulCtrlMP.scala 170:30]
      uart_buffer <= 8'h0; // @[NulCtrlMP.scala 170:30]
    end else if (state == 5'h19) begin // @[NulCtrlMP.scala 938:29]
      if (send_hear) begin // @[NulCtrlMP.scala 939:20]
        if (_T_672) begin // @[NulCtrlMP.scala 943:23]
          uart_buffer <= 8'h0; // @[NulCtrlMP.scala 945:21]
        end
      end else if (_T_674) begin // @[NulCtrlMP.scala 953:23]
        uart_buffer <= io_rx_bits; // @[NulCtrlMP.scala 954:21]
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 172:28]
      sleep_cnt <= 4'h0; // @[NulCtrlMP.scala 172:28]
    end else if (state == 5'h1f) begin // @[NulCtrlMP.scala 173:33]
      sleep_cnt <= _sleep_cnt_T_1; // @[NulCtrlMP.scala 174:19]
    end
    cnt <= _GEN_10151[127:0]; // @[NulCtrlMP.scala 345:{22,22}]
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_0 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[0]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_0 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end else begin
          regback_0 <= _GEN_7348;
        end
      end else begin
        regback_0 <= _GEN_7348;
      end
    end else begin
      regback_0 <= _GEN_7348;
    end
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_1 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[1]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_1 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end else begin
          regback_1 <= _GEN_7349;
        end
      end else begin
        regback_1 <= _GEN_7349;
      end
    end else begin
      regback_1 <= _GEN_7349;
    end
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_2 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[2]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_2 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end else begin
          regback_2 <= _GEN_7350;
        end
      end else begin
        regback_2 <= _GEN_7350;
      end
    end else begin
      regback_2 <= _GEN_7350;
    end
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_3 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[3]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_3 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end else begin
          regback_3 <= _GEN_7351;
        end
      end else begin
        regback_3 <= _GEN_7351;
      end
    end else begin
      regback_3 <= _GEN_7351;
    end
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_4 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[4]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_4 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end else begin
          regback_4 <= _GEN_7352;
        end
      end else begin
        regback_4 <= _GEN_7352;
      end
    end else begin
      regback_4 <= _GEN_7352;
    end
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_5 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[5]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_5 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end else begin
          regback_5 <= _GEN_7353;
        end
      end else begin
        regback_5 <= _GEN_7353;
      end
    end else begin
      regback_5 <= _GEN_7353;
    end
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_6 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[6]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_6 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end else begin
          regback_6 <= _GEN_7354;
        end
      end else begin
        regback_6 <= _GEN_7354;
      end
    end else begin
      regback_6 <= _GEN_7354;
    end
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_7 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[7]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_7 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end else begin
          regback_7 <= _GEN_7355;
        end
      end else begin
        regback_7 <= _GEN_7355;
      end
    end else begin
      regback_7 <= _GEN_7355;
    end
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_8 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[8]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_8 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end else begin
          regback_8 <= _GEN_7356;
        end
      end else begin
        regback_8 <= _GEN_7356;
      end
    end else begin
      regback_8 <= _GEN_7356;
    end
    if (reset) begin // @[NulCtrlMP.scala 346:26]
      regback_9 <= 64'h0; // @[NulCtrlMP.scala 346:26]
    end else if (state == 5'h15) begin // @[NulCtrlMP.scala 777:32]
      if (cnt[9]) begin // @[NulCtrlMP.scala 408:32]
        if (_T_122) begin // @[NulCtrlMP.scala 353:36]
          regback_9 <= _GEN_1349; // @[NulCtrlMP.scala 355:17]
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 420:27]
      init_cnt <= 2'h0; // @[NulCtrlMP.scala 420:27]
    end else if (state == 5'h1) begin // @[NulCtrlMP.scala 421:35]
      if (cnt[8]) begin // @[NulCtrlMP.scala 442:22]
        if (!(init_cnt == 2'h3)) begin // @[NulCtrlMP.scala 444:47]
          init_cnt <= _nextidx_T_1; // @[NulCtrlMP.scala 449:26]
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 742:30]
      pg_loop_cnt <= 8'h0; // @[NulCtrlMP.scala 742:30]
    end else if (state == 5'h15) begin // @[NulCtrlMP.scala 777:32]
      if (cnt[31]) begin // @[NulCtrlMP.scala 800:23]
        if (pg_loop_cnt < 8'h3f) begin // @[NulCtrlMP.scala 801:38]
          pg_loop_cnt <= _pg_loop_cnt_T_1; // @[NulCtrlMP.scala 803:29]
        end else begin
          pg_loop_cnt <= 8'h0; // @[NulCtrlMP.scala 806:29]
        end
      end else begin
        pg_loop_cnt <= _GEN_4013;
      end
    end else begin
      pg_loop_cnt <= _GEN_4013;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_0 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_0 <= _GEN_7455;
        end else begin
          pgbuf_div8_0 <= _GEN_7379;
        end
      end else begin
        pgbuf_div8_0 <= _GEN_7379;
      end
    end else begin
      pgbuf_div8_0 <= _GEN_7379;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_1 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_1 <= _GEN_7456;
        end else begin
          pgbuf_div8_1 <= _GEN_7380;
        end
      end else begin
        pgbuf_div8_1 <= _GEN_7380;
      end
    end else begin
      pgbuf_div8_1 <= _GEN_7380;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_2 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_2 <= _GEN_7457;
        end else begin
          pgbuf_div8_2 <= _GEN_7381;
        end
      end else begin
        pgbuf_div8_2 <= _GEN_7381;
      end
    end else begin
      pgbuf_div8_2 <= _GEN_7381;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_3 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_3 <= _GEN_7458;
        end else begin
          pgbuf_div8_3 <= _GEN_7382;
        end
      end else begin
        pgbuf_div8_3 <= _GEN_7382;
      end
    end else begin
      pgbuf_div8_3 <= _GEN_7382;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_4 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_4 <= _GEN_7459;
        end else begin
          pgbuf_div8_4 <= _GEN_7383;
        end
      end else begin
        pgbuf_div8_4 <= _GEN_7383;
      end
    end else begin
      pgbuf_div8_4 <= _GEN_7383;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_5 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_5 <= _GEN_7460;
        end else begin
          pgbuf_div8_5 <= _GEN_7384;
        end
      end else begin
        pgbuf_div8_5 <= _GEN_7384;
      end
    end else begin
      pgbuf_div8_5 <= _GEN_7384;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_6 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_6 <= _GEN_7461;
        end else begin
          pgbuf_div8_6 <= _GEN_7385;
        end
      end else begin
        pgbuf_div8_6 <= _GEN_7385;
      end
    end else begin
      pgbuf_div8_6 <= _GEN_7385;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_7 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_7 <= _GEN_7462;
        end else begin
          pgbuf_div8_7 <= _GEN_7386;
        end
      end else begin
        pgbuf_div8_7 <= _GEN_7386;
      end
    end else begin
      pgbuf_div8_7 <= _GEN_7386;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_8 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_8 <= _GEN_7463;
        end else begin
          pgbuf_div8_8 <= _GEN_7387;
        end
      end else begin
        pgbuf_div8_8 <= _GEN_7387;
      end
    end else begin
      pgbuf_div8_8 <= _GEN_7387;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_9 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_9 <= _GEN_7464;
        end else begin
          pgbuf_div8_9 <= _GEN_7388;
        end
      end else begin
        pgbuf_div8_9 <= _GEN_7388;
      end
    end else begin
      pgbuf_div8_9 <= _GEN_7388;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_10 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_10 <= _GEN_7465;
        end else begin
          pgbuf_div8_10 <= _GEN_7389;
        end
      end else begin
        pgbuf_div8_10 <= _GEN_7389;
      end
    end else begin
      pgbuf_div8_10 <= _GEN_7389;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_11 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_11 <= _GEN_7466;
        end else begin
          pgbuf_div8_11 <= _GEN_7390;
        end
      end else begin
        pgbuf_div8_11 <= _GEN_7390;
      end
    end else begin
      pgbuf_div8_11 <= _GEN_7390;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_12 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_12 <= _GEN_7467;
        end else begin
          pgbuf_div8_12 <= _GEN_7391;
        end
      end else begin
        pgbuf_div8_12 <= _GEN_7391;
      end
    end else begin
      pgbuf_div8_12 <= _GEN_7391;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_13 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_13 <= _GEN_7468;
        end else begin
          pgbuf_div8_13 <= _GEN_7392;
        end
      end else begin
        pgbuf_div8_13 <= _GEN_7392;
      end
    end else begin
      pgbuf_div8_13 <= _GEN_7392;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_14 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_14 <= _GEN_7469;
        end else begin
          pgbuf_div8_14 <= _GEN_7393;
        end
      end else begin
        pgbuf_div8_14 <= _GEN_7393;
      end
    end else begin
      pgbuf_div8_14 <= _GEN_7393;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_15 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_15 <= _GEN_7470;
        end else begin
          pgbuf_div8_15 <= _GEN_7394;
        end
      end else begin
        pgbuf_div8_15 <= _GEN_7394;
      end
    end else begin
      pgbuf_div8_15 <= _GEN_7394;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_16 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_16 <= _GEN_7471;
        end else begin
          pgbuf_div8_16 <= _GEN_7395;
        end
      end else begin
        pgbuf_div8_16 <= _GEN_7395;
      end
    end else begin
      pgbuf_div8_16 <= _GEN_7395;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_17 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_17 <= _GEN_7472;
        end else begin
          pgbuf_div8_17 <= _GEN_7396;
        end
      end else begin
        pgbuf_div8_17 <= _GEN_7396;
      end
    end else begin
      pgbuf_div8_17 <= _GEN_7396;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_18 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_18 <= _GEN_7473;
        end else begin
          pgbuf_div8_18 <= _GEN_7397;
        end
      end else begin
        pgbuf_div8_18 <= _GEN_7397;
      end
    end else begin
      pgbuf_div8_18 <= _GEN_7397;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_19 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_19 <= _GEN_7474;
        end else begin
          pgbuf_div8_19 <= _GEN_7398;
        end
      end else begin
        pgbuf_div8_19 <= _GEN_7398;
      end
    end else begin
      pgbuf_div8_19 <= _GEN_7398;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_20 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_20 <= _GEN_7475;
        end else begin
          pgbuf_div8_20 <= _GEN_7399;
        end
      end else begin
        pgbuf_div8_20 <= _GEN_7399;
      end
    end else begin
      pgbuf_div8_20 <= _GEN_7399;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_21 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_21 <= _GEN_7476;
        end else begin
          pgbuf_div8_21 <= _GEN_7400;
        end
      end else begin
        pgbuf_div8_21 <= _GEN_7400;
      end
    end else begin
      pgbuf_div8_21 <= _GEN_7400;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_22 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_22 <= _GEN_7477;
        end else begin
          pgbuf_div8_22 <= _GEN_7401;
        end
      end else begin
        pgbuf_div8_22 <= _GEN_7401;
      end
    end else begin
      pgbuf_div8_22 <= _GEN_7401;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_23 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_23 <= _GEN_7478;
        end else begin
          pgbuf_div8_23 <= _GEN_7402;
        end
      end else begin
        pgbuf_div8_23 <= _GEN_7402;
      end
    end else begin
      pgbuf_div8_23 <= _GEN_7402;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_24 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_24 <= _GEN_7479;
        end else begin
          pgbuf_div8_24 <= _GEN_7403;
        end
      end else begin
        pgbuf_div8_24 <= _GEN_7403;
      end
    end else begin
      pgbuf_div8_24 <= _GEN_7403;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_25 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_25 <= _GEN_7480;
        end else begin
          pgbuf_div8_25 <= _GEN_7404;
        end
      end else begin
        pgbuf_div8_25 <= _GEN_7404;
      end
    end else begin
      pgbuf_div8_25 <= _GEN_7404;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_26 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_26 <= _GEN_7481;
        end else begin
          pgbuf_div8_26 <= _GEN_7405;
        end
      end else begin
        pgbuf_div8_26 <= _GEN_7405;
      end
    end else begin
      pgbuf_div8_26 <= _GEN_7405;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_27 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_27 <= _GEN_7482;
        end else begin
          pgbuf_div8_27 <= _GEN_7406;
        end
      end else begin
        pgbuf_div8_27 <= _GEN_7406;
      end
    end else begin
      pgbuf_div8_27 <= _GEN_7406;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_28 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_28 <= _GEN_7483;
        end else begin
          pgbuf_div8_28 <= _GEN_7407;
        end
      end else begin
        pgbuf_div8_28 <= _GEN_7407;
      end
    end else begin
      pgbuf_div8_28 <= _GEN_7407;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_29 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_29 <= _GEN_7484;
        end else begin
          pgbuf_div8_29 <= _GEN_7408;
        end
      end else begin
        pgbuf_div8_29 <= _GEN_7408;
      end
    end else begin
      pgbuf_div8_29 <= _GEN_7408;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_30 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_30 <= _GEN_7485;
        end else begin
          pgbuf_div8_30 <= _GEN_7409;
        end
      end else begin
        pgbuf_div8_30 <= _GEN_7409;
      end
    end else begin
      pgbuf_div8_30 <= _GEN_7409;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_31 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_31 <= _GEN_7486;
        end else begin
          pgbuf_div8_31 <= _GEN_7410;
        end
      end else begin
        pgbuf_div8_31 <= _GEN_7410;
      end
    end else begin
      pgbuf_div8_31 <= _GEN_7410;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_32 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_32 <= _GEN_7487;
        end else begin
          pgbuf_div8_32 <= _GEN_7411;
        end
      end else begin
        pgbuf_div8_32 <= _GEN_7411;
      end
    end else begin
      pgbuf_div8_32 <= _GEN_7411;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_33 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_33 <= _GEN_7488;
        end else begin
          pgbuf_div8_33 <= _GEN_7412;
        end
      end else begin
        pgbuf_div8_33 <= _GEN_7412;
      end
    end else begin
      pgbuf_div8_33 <= _GEN_7412;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_34 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_34 <= _GEN_7489;
        end else begin
          pgbuf_div8_34 <= _GEN_7413;
        end
      end else begin
        pgbuf_div8_34 <= _GEN_7413;
      end
    end else begin
      pgbuf_div8_34 <= _GEN_7413;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_35 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_35 <= _GEN_7490;
        end else begin
          pgbuf_div8_35 <= _GEN_7414;
        end
      end else begin
        pgbuf_div8_35 <= _GEN_7414;
      end
    end else begin
      pgbuf_div8_35 <= _GEN_7414;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_36 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_36 <= _GEN_7491;
        end else begin
          pgbuf_div8_36 <= _GEN_7415;
        end
      end else begin
        pgbuf_div8_36 <= _GEN_7415;
      end
    end else begin
      pgbuf_div8_36 <= _GEN_7415;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_37 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_37 <= _GEN_7492;
        end else begin
          pgbuf_div8_37 <= _GEN_7416;
        end
      end else begin
        pgbuf_div8_37 <= _GEN_7416;
      end
    end else begin
      pgbuf_div8_37 <= _GEN_7416;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_38 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_38 <= _GEN_7493;
        end else begin
          pgbuf_div8_38 <= _GEN_7417;
        end
      end else begin
        pgbuf_div8_38 <= _GEN_7417;
      end
    end else begin
      pgbuf_div8_38 <= _GEN_7417;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_39 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_39 <= _GEN_7494;
        end else begin
          pgbuf_div8_39 <= _GEN_7418;
        end
      end else begin
        pgbuf_div8_39 <= _GEN_7418;
      end
    end else begin
      pgbuf_div8_39 <= _GEN_7418;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_40 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_40 <= _GEN_7495;
        end else begin
          pgbuf_div8_40 <= _GEN_7419;
        end
      end else begin
        pgbuf_div8_40 <= _GEN_7419;
      end
    end else begin
      pgbuf_div8_40 <= _GEN_7419;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_41 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_41 <= _GEN_7496;
        end else begin
          pgbuf_div8_41 <= _GEN_7420;
        end
      end else begin
        pgbuf_div8_41 <= _GEN_7420;
      end
    end else begin
      pgbuf_div8_41 <= _GEN_7420;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_42 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_42 <= _GEN_7497;
        end else begin
          pgbuf_div8_42 <= _GEN_7421;
        end
      end else begin
        pgbuf_div8_42 <= _GEN_7421;
      end
    end else begin
      pgbuf_div8_42 <= _GEN_7421;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_43 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_43 <= _GEN_7498;
        end else begin
          pgbuf_div8_43 <= _GEN_7422;
        end
      end else begin
        pgbuf_div8_43 <= _GEN_7422;
      end
    end else begin
      pgbuf_div8_43 <= _GEN_7422;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_44 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_44 <= _GEN_7499;
        end else begin
          pgbuf_div8_44 <= _GEN_7423;
        end
      end else begin
        pgbuf_div8_44 <= _GEN_7423;
      end
    end else begin
      pgbuf_div8_44 <= _GEN_7423;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_45 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_45 <= _GEN_7500;
        end else begin
          pgbuf_div8_45 <= _GEN_7424;
        end
      end else begin
        pgbuf_div8_45 <= _GEN_7424;
      end
    end else begin
      pgbuf_div8_45 <= _GEN_7424;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_46 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_46 <= _GEN_7501;
        end else begin
          pgbuf_div8_46 <= _GEN_7425;
        end
      end else begin
        pgbuf_div8_46 <= _GEN_7425;
      end
    end else begin
      pgbuf_div8_46 <= _GEN_7425;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_47 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_47 <= _GEN_7502;
        end else begin
          pgbuf_div8_47 <= _GEN_7426;
        end
      end else begin
        pgbuf_div8_47 <= _GEN_7426;
      end
    end else begin
      pgbuf_div8_47 <= _GEN_7426;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_48 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_48 <= _GEN_7503;
        end else begin
          pgbuf_div8_48 <= _GEN_7427;
        end
      end else begin
        pgbuf_div8_48 <= _GEN_7427;
      end
    end else begin
      pgbuf_div8_48 <= _GEN_7427;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_49 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_49 <= _GEN_7504;
        end else begin
          pgbuf_div8_49 <= _GEN_7428;
        end
      end else begin
        pgbuf_div8_49 <= _GEN_7428;
      end
    end else begin
      pgbuf_div8_49 <= _GEN_7428;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_50 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_50 <= _GEN_7505;
        end else begin
          pgbuf_div8_50 <= _GEN_7429;
        end
      end else begin
        pgbuf_div8_50 <= _GEN_7429;
      end
    end else begin
      pgbuf_div8_50 <= _GEN_7429;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_51 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_51 <= _GEN_7506;
        end else begin
          pgbuf_div8_51 <= _GEN_7430;
        end
      end else begin
        pgbuf_div8_51 <= _GEN_7430;
      end
    end else begin
      pgbuf_div8_51 <= _GEN_7430;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_52 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_52 <= _GEN_7507;
        end else begin
          pgbuf_div8_52 <= _GEN_7431;
        end
      end else begin
        pgbuf_div8_52 <= _GEN_7431;
      end
    end else begin
      pgbuf_div8_52 <= _GEN_7431;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_53 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_53 <= _GEN_7508;
        end else begin
          pgbuf_div8_53 <= _GEN_7432;
        end
      end else begin
        pgbuf_div8_53 <= _GEN_7432;
      end
    end else begin
      pgbuf_div8_53 <= _GEN_7432;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_54 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_54 <= _GEN_7509;
        end else begin
          pgbuf_div8_54 <= _GEN_7433;
        end
      end else begin
        pgbuf_div8_54 <= _GEN_7433;
      end
    end else begin
      pgbuf_div8_54 <= _GEN_7433;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_55 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_55 <= _GEN_7510;
        end else begin
          pgbuf_div8_55 <= _GEN_7434;
        end
      end else begin
        pgbuf_div8_55 <= _GEN_7434;
      end
    end else begin
      pgbuf_div8_55 <= _GEN_7434;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_56 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_56 <= _GEN_7511;
        end else begin
          pgbuf_div8_56 <= _GEN_7435;
        end
      end else begin
        pgbuf_div8_56 <= _GEN_7435;
      end
    end else begin
      pgbuf_div8_56 <= _GEN_7435;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_57 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_57 <= _GEN_7512;
        end else begin
          pgbuf_div8_57 <= _GEN_7436;
        end
      end else begin
        pgbuf_div8_57 <= _GEN_7436;
      end
    end else begin
      pgbuf_div8_57 <= _GEN_7436;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_58 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_58 <= _GEN_7513;
        end else begin
          pgbuf_div8_58 <= _GEN_7437;
        end
      end else begin
        pgbuf_div8_58 <= _GEN_7437;
      end
    end else begin
      pgbuf_div8_58 <= _GEN_7437;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_59 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_59 <= _GEN_7514;
        end else begin
          pgbuf_div8_59 <= _GEN_7438;
        end
      end else begin
        pgbuf_div8_59 <= _GEN_7438;
      end
    end else begin
      pgbuf_div8_59 <= _GEN_7438;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_60 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_60 <= _GEN_7515;
        end else begin
          pgbuf_div8_60 <= _GEN_7439;
        end
      end else begin
        pgbuf_div8_60 <= _GEN_7439;
      end
    end else begin
      pgbuf_div8_60 <= _GEN_7439;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_61 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_61 <= _GEN_7516;
        end else begin
          pgbuf_div8_61 <= _GEN_7440;
        end
      end else begin
        pgbuf_div8_61 <= _GEN_7440;
      end
    end else begin
      pgbuf_div8_61 <= _GEN_7440;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_62 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_62 <= _GEN_7517;
        end else begin
          pgbuf_div8_62 <= _GEN_7441;
        end
      end else begin
        pgbuf_div8_62 <= _GEN_7441;
      end
    end else begin
      pgbuf_div8_62 <= _GEN_7441;
    end
    if (reset) begin // @[NulCtrlMP.scala 818:29]
      pgbuf_div8_63 <= 64'h0; // @[NulCtrlMP.scala 818:29]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (wt_byte_cnt == 4'h7) begin // @[NulCtrlMP.scala 885:39]
          pgbuf_div8_63 <= _GEN_7518;
        end else begin
          pgbuf_div8_63 <= _GEN_7442;
        end
      end else begin
        pgbuf_div8_63 <= _GEN_7442;
      end
    end else begin
      pgbuf_div8_63 <= _GEN_7442;
    end
    if (reset) begin // @[NulCtrlMP.scala 819:33]
      pgbuf_uart_pos <= 12'h0; // @[NulCtrlMP.scala 819:33]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[41]) begin // @[NulCtrlMP.scala 925:23]
        pgbuf_uart_pos <= 12'h0; // @[NulCtrlMP.scala 929:28]
      end else if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        pgbuf_uart_pos <= _GEN_7584;
      end else begin
        pgbuf_uart_pos <= _GEN_7445;
      end
    end else begin
      pgbuf_uart_pos <= _GEN_7445;
    end
    if (reset) begin // @[NulCtrlMP.scala 820:32]
      pgbuf_cpu_pos <= 12'h0; // @[NulCtrlMP.scala 820:32]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[41]) begin // @[NulCtrlMP.scala 925:23]
        pgbuf_cpu_pos <= 12'h0; // @[NulCtrlMP.scala 928:27]
      end else if (cnt[29]) begin // @[NulCtrlMP.scala 914:23]
        pgbuf_cpu_pos <= _pgbuf_cpu_pos_T_1; // @[NulCtrlMP.scala 920:27]
      end else begin
        pgbuf_cpu_pos <= _GEN_7443;
      end
    end else begin
      pgbuf_cpu_pos <= _GEN_7443;
    end
    if (reset) begin // @[NulCtrlMP.scala 876:30]
      wt_byte_cnt <= 4'h0; // @[NulCtrlMP.scala 876:30]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (cnt[41]) begin // @[NulCtrlMP.scala 925:23]
        wt_byte_cnt <= 4'h0; // @[NulCtrlMP.scala 930:25]
      end else if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        wt_byte_cnt <= _GEN_7519;
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 877:30]
      wt_byte_buf_0 <= 8'h0; // @[NulCtrlMP.scala 877:30]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (3'h0 == wt_byte_cnt[2:0]) begin // @[NulCtrlMP.scala 884:38]
          wt_byte_buf_0 <= io_rx_bits; // @[NulCtrlMP.scala 884:38]
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 877:30]
      wt_byte_buf_1 <= 8'h0; // @[NulCtrlMP.scala 877:30]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (3'h1 == wt_byte_cnt[2:0]) begin // @[NulCtrlMP.scala 884:38]
          wt_byte_buf_1 <= io_rx_bits; // @[NulCtrlMP.scala 884:38]
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 877:30]
      wt_byte_buf_2 <= 8'h0; // @[NulCtrlMP.scala 877:30]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (3'h2 == wt_byte_cnt[2:0]) begin // @[NulCtrlMP.scala 884:38]
          wt_byte_buf_2 <= io_rx_bits; // @[NulCtrlMP.scala 884:38]
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 877:30]
      wt_byte_buf_3 <= 8'h0; // @[NulCtrlMP.scala 877:30]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (3'h3 == wt_byte_cnt[2:0]) begin // @[NulCtrlMP.scala 884:38]
          wt_byte_buf_3 <= io_rx_bits; // @[NulCtrlMP.scala 884:38]
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 877:30]
      wt_byte_buf_4 <= 8'h0; // @[NulCtrlMP.scala 877:30]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (3'h4 == wt_byte_cnt[2:0]) begin // @[NulCtrlMP.scala 884:38]
          wt_byte_buf_4 <= io_rx_bits; // @[NulCtrlMP.scala 884:38]
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 877:30]
      wt_byte_buf_5 <= 8'h0; // @[NulCtrlMP.scala 877:30]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (3'h5 == wt_byte_cnt[2:0]) begin // @[NulCtrlMP.scala 884:38]
          wt_byte_buf_5 <= io_rx_bits; // @[NulCtrlMP.scala 884:38]
        end
      end
    end
    if (reset) begin // @[NulCtrlMP.scala 877:30]
      wt_byte_buf_6 <= 8'h0; // @[NulCtrlMP.scala 877:30]
    end else if (state == 5'h14) begin // @[NulCtrlMP.scala 879:32]
      if (io_rx_valid & _T_555) begin // @[NulCtrlMP.scala 883:55]
        if (3'h6 == wt_byte_cnt[2:0]) begin // @[NulCtrlMP.scala 884:38]
          wt_byte_buf_6 <= io_rx_bits; // @[NulCtrlMP.scala 884:38]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cpu_state_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_state_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  cpu_state_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  cpu_state_3 = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  global_clk = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  user_clk_0 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  user_clk_1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  user_clk_2 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  user_clk_3 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  cpu_raised_itr_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  cpu_raised_itr_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cpu_raised_itr_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  cpu_raised_itr_3 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  last_priv_0 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  last_priv_1 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  last_priv_2 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  last_priv_3 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  state = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  trans_bytes = _RAND_18[9:0];
  _RAND_19 = {1{`RANDOM}};
  trans_pos = _RAND_19[9:0];
  _RAND_20 = {1{`RANDOM}};
  errno = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  opcode = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  opoff = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  oparg_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  oparg_2 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  oparg_3 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  oparg_4 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  oparg_5 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  oparg_6 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  oparg_7 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  oparg_8 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  oparg_9 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  oparg_10 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  oparg_11 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  oparg_12 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  oparg_13 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  oparg_14 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  oparg_15 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  retarg_0 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  retarg_1 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  retarg_2 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  retarg_3 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  retarg_4 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  retarg_5 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  retarg_6 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  retarg_7 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  retarg_8 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  retarg_9 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  retarg_10 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  retarg_11 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  retarg_12 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  retarg_13 = _RAND_51[7:0];
  _RAND_52 = {2{`RANDOM}};
  hfutex_masks_0_0 = _RAND_52[47:0];
  _RAND_53 = {2{`RANDOM}};
  hfutex_masks_0_1 = _RAND_53[47:0];
  _RAND_54 = {2{`RANDOM}};
  hfutex_masks_0_2 = _RAND_54[47:0];
  _RAND_55 = {2{`RANDOM}};
  hfutex_masks_0_3 = _RAND_55[47:0];
  _RAND_56 = {2{`RANDOM}};
  hfutex_masks_1_0 = _RAND_56[47:0];
  _RAND_57 = {2{`RANDOM}};
  hfutex_masks_1_1 = _RAND_57[47:0];
  _RAND_58 = {2{`RANDOM}};
  hfutex_masks_1_2 = _RAND_58[47:0];
  _RAND_59 = {2{`RANDOM}};
  hfutex_masks_1_3 = _RAND_59[47:0];
  _RAND_60 = {2{`RANDOM}};
  hfutex_masks_2_0 = _RAND_60[47:0];
  _RAND_61 = {2{`RANDOM}};
  hfutex_masks_2_1 = _RAND_61[47:0];
  _RAND_62 = {2{`RANDOM}};
  hfutex_masks_2_2 = _RAND_62[47:0];
  _RAND_63 = {2{`RANDOM}};
  hfutex_masks_2_3 = _RAND_63[47:0];
  _RAND_64 = {2{`RANDOM}};
  hfutex_masks_3_0 = _RAND_64[47:0];
  _RAND_65 = {2{`RANDOM}};
  hfutex_masks_3_1 = _RAND_65[47:0];
  _RAND_66 = {2{`RANDOM}};
  hfutex_masks_3_2 = _RAND_66[47:0];
  _RAND_67 = {2{`RANDOM}};
  hfutex_masks_3_3 = _RAND_67[47:0];
  _RAND_68 = {1{`RANDOM}};
  hfutex_pos_0 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  hfutex_pos_1 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  hfutex_pos_2 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  hfutex_pos_3 = _RAND_71[1:0];
  _RAND_72 = {2{`RANDOM}};
  hfutex_match_reg = _RAND_72[47:0];
  _RAND_73 = {1{`RANDOM}};
  send_hear = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  uart_buffer = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  sleep_cnt = _RAND_75[3:0];
  _RAND_76 = {4{`RANDOM}};
  cnt = _RAND_76[127:0];
  _RAND_77 = {2{`RANDOM}};
  regback_0 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  regback_1 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  regback_2 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  regback_3 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  regback_4 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  regback_5 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  regback_6 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  regback_7 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  regback_8 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  regback_9 = _RAND_86[63:0];
  _RAND_87 = {1{`RANDOM}};
  init_cnt = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  pg_loop_cnt = _RAND_88[7:0];
  _RAND_89 = {2{`RANDOM}};
  pgbuf_div8_0 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  pgbuf_div8_1 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  pgbuf_div8_2 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  pgbuf_div8_3 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  pgbuf_div8_4 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  pgbuf_div8_5 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  pgbuf_div8_6 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  pgbuf_div8_7 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  pgbuf_div8_8 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  pgbuf_div8_9 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  pgbuf_div8_10 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  pgbuf_div8_11 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  pgbuf_div8_12 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  pgbuf_div8_13 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  pgbuf_div8_14 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  pgbuf_div8_15 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  pgbuf_div8_16 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  pgbuf_div8_17 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  pgbuf_div8_18 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  pgbuf_div8_19 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  pgbuf_div8_20 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  pgbuf_div8_21 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  pgbuf_div8_22 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  pgbuf_div8_23 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  pgbuf_div8_24 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  pgbuf_div8_25 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  pgbuf_div8_26 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  pgbuf_div8_27 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  pgbuf_div8_28 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  pgbuf_div8_29 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  pgbuf_div8_30 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  pgbuf_div8_31 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  pgbuf_div8_32 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  pgbuf_div8_33 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  pgbuf_div8_34 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  pgbuf_div8_35 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  pgbuf_div8_36 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  pgbuf_div8_37 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  pgbuf_div8_38 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  pgbuf_div8_39 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  pgbuf_div8_40 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  pgbuf_div8_41 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  pgbuf_div8_42 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  pgbuf_div8_43 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  pgbuf_div8_44 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  pgbuf_div8_45 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  pgbuf_div8_46 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  pgbuf_div8_47 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  pgbuf_div8_48 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  pgbuf_div8_49 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  pgbuf_div8_50 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  pgbuf_div8_51 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  pgbuf_div8_52 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  pgbuf_div8_53 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  pgbuf_div8_54 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  pgbuf_div8_55 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  pgbuf_div8_56 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  pgbuf_div8_57 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  pgbuf_div8_58 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  pgbuf_div8_59 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  pgbuf_div8_60 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  pgbuf_div8_61 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  pgbuf_div8_62 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  pgbuf_div8_63 = _RAND_152[63:0];
  _RAND_153 = {1{`RANDOM}};
  pgbuf_uart_pos = _RAND_153[11:0];
  _RAND_154 = {1{`RANDOM}};
  pgbuf_cpu_pos = _RAND_154[11:0];
  _RAND_155 = {1{`RANDOM}};
  wt_byte_cnt = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  wt_byte_buf_0 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  wt_byte_buf_1 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  wt_byte_buf_2 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  wt_byte_buf_3 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  wt_byte_buf_4 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  wt_byte_buf_5 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  wt_byte_buf_6 = _RAND_162[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Tx(
  input        clock,
  input        reset,
  output       io_txd,
  output       io_channel_ready,
  input        io_channel_valid,
  input  [7:0] io_channel_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [10:0] shiftReg; // @[port.scala 39:27]
  reg [19:0] cntReg; // @[port.scala 40:25]
  reg [3:0] bitsReg; // @[port.scala 41:26]
  wire  _io_channel_ready_T = cntReg == 20'h0; // @[port.scala 43:33]
  wire [9:0] shift = shiftReg[10:1]; // @[port.scala 50:34]
  wire [10:0] _shiftReg_T_1 = {1'h1,shift}; // @[port.scala 51:29]
  wire [3:0] _bitsReg_T_1 = bitsReg - 4'h1; // @[port.scala 52:32]
  wire [10:0] _shiftReg_T_3 = {2'h3,io_channel_bits,1'h0}; // @[port.scala 56:52]
  wire [19:0] _cntReg_T_1 = cntReg - 20'h1; // @[port.scala 64:26]
  assign io_txd = shiftReg[0]; // @[port.scala 44:23]
  assign io_channel_ready = cntReg == 20'h0 & bitsReg == 4'h0; // @[port.scala 43:42]
  always @(posedge clock) begin
    if (reset) begin // @[port.scala 39:27]
      shiftReg <= 11'h7ff; // @[port.scala 39:27]
    end else if (_io_channel_ready_T) begin // @[port.scala 46:26]
      if (bitsReg != 4'h0) begin // @[port.scala 49:31]
        shiftReg <= _shiftReg_T_1; // @[port.scala 51:22]
      end else if (io_channel_valid) begin // @[port.scala 54:36]
        shiftReg <= _shiftReg_T_3; // @[port.scala 56:26]
      end else begin
        shiftReg <= 11'h7ff; // @[port.scala 59:26]
      end
    end
    if (reset) begin // @[port.scala 40:25]
      cntReg <= 20'h0; // @[port.scala 40:25]
    end else if (_io_channel_ready_T) begin // @[port.scala 46:26]
      cntReg <= 20'h6c; // @[port.scala 48:16]
    end else begin
      cntReg <= _cntReg_T_1; // @[port.scala 64:16]
    end
    if (reset) begin // @[port.scala 41:26]
      bitsReg <= 4'h0; // @[port.scala 41:26]
    end else if (_io_channel_ready_T) begin // @[port.scala 46:26]
      if (bitsReg != 4'h0) begin // @[port.scala 49:31]
        bitsReg <= _bitsReg_T_1; // @[port.scala 52:21]
      end else if (io_channel_valid) begin // @[port.scala 54:36]
        bitsReg <= 4'hb; // @[port.scala 57:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shiftReg = _RAND_0[10:0];
  _RAND_1 = {1{`RANDOM}};
  cntReg = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  bitsReg = _RAND_2[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Rx(
  input        clock,
  input        reset,
  input        io_rxd,
  input        io_channel_ready,
  output       io_channel_valid,
  output [7:0] io_channel_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  rxReg_REG; // @[port.scala 80:32]
  reg  rxReg; // @[port.scala 80:24]
  reg [7:0] shiftReg; // @[port.scala 82:27]
  reg [19:0] cntReg; // @[port.scala 83:25]
  reg [3:0] bitsReg; // @[port.scala 84:26]
  reg  validReg; // @[port.scala 85:27]
  wire [19:0] _cntReg_T_1 = cntReg - 20'h1; // @[port.scala 88:26]
  wire [7:0] _shiftReg_T_1 = {rxReg,shiftReg[7:1]}; // @[port.scala 91:27]
  wire [3:0] _bitsReg_T_1 = bitsReg - 4'h1; // @[port.scala 92:28]
  wire  _GEN_0 = bitsReg == 4'h1 | validReg; // @[port.scala 94:31 95:18 85:27]
  assign io_channel_valid = validReg; // @[port.scala 108:22]
  assign io_channel_bits = shiftReg; // @[port.scala 107:21]
  always @(posedge clock) begin
    rxReg_REG <= reset | io_rxd; // @[port.scala 80:{32,32,32}]
    rxReg <= reset | rxReg_REG; // @[port.scala 80:{24,24,24}]
    if (reset) begin // @[port.scala 82:27]
      shiftReg <= 8'h0; // @[port.scala 82:27]
    end else if (!(cntReg != 20'h0)) begin // @[port.scala 87:26]
      if (bitsReg != 4'h0) begin // @[port.scala 89:34]
        shiftReg <= _shiftReg_T_1; // @[port.scala 91:18]
      end
    end
    if (reset) begin // @[port.scala 83:25]
      cntReg <= 20'h0; // @[port.scala 83:25]
    end else if (cntReg != 20'h0) begin // @[port.scala 87:26]
      cntReg <= _cntReg_T_1; // @[port.scala 88:16]
    end else if (bitsReg != 4'h0) begin // @[port.scala 89:34]
      cntReg <= 20'h6c; // @[port.scala 90:16]
    end else if (~rxReg) begin // @[port.scala 97:32]
      cntReg <= 20'ha2; // @[port.scala 99:16]
    end
    if (reset) begin // @[port.scala 84:26]
      bitsReg <= 4'h0; // @[port.scala 84:26]
    end else if (!(cntReg != 20'h0)) begin // @[port.scala 87:26]
      if (bitsReg != 4'h0) begin // @[port.scala 89:34]
        bitsReg <= _bitsReg_T_1; // @[port.scala 92:17]
      end else if (~rxReg) begin // @[port.scala 97:32]
        bitsReg <= 4'h8; // @[port.scala 100:17]
      end
    end
    if (reset) begin // @[port.scala 85:27]
      validReg <= 1'h0; // @[port.scala 85:27]
    end else if (validReg & io_channel_ready) begin // @[port.scala 103:40]
      validReg <= 1'h0; // @[port.scala 104:18]
    end else if (!(cntReg != 20'h0)) begin // @[port.scala 87:26]
      if (bitsReg != 4'h0) begin // @[port.scala 89:34]
        validReg <= _GEN_0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rxReg_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  rxReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shiftReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  cntReg = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  bitsReg = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  validReg = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output [9:0] io_count
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:511]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [8:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire [8:0] ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg [8:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [8:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [8:0] _value_T_1 = enq_ptr_value + 9'h1; // @[Counter.scala 78:24]
  wire [8:0] _value_T_3 = deq_ptr_value + 9'h1; // @[Counter.scala 78:24]
  wire [8:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 312:32]
  wire [9:0] _io_count_T_1 = maybe_full & ptr_match ? 10'h200 : 10'h0; // @[Decoupled.scala 315:20]
  wire [9:0] _GEN_11 = {{1'd0}, ptr_diff}; // @[Decoupled.scala 315:62]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_count = _io_count_T_1 | _GEN_11; // @[Decoupled.scala 315:62]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 9'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 9'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_2(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [5:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _value_T_1 = enq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire [5:0] _value_T_3 = deq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NulCPUCtrlMPWithUart(
  input         clock,
  input         reset,
  input         io_cpu_0_inited,
  input  [1:0]  io_cpu_0_priv,
  output        io_cpu_0_ext_itr,
  output        io_cpu_0_stop_fetch,
  output        io_cpu_0_regacc_rd,
  output        io_cpu_0_regacc_wt,
  output [4:0]  io_cpu_0_regacc_idx,
  output [63:0] io_cpu_0_regacc_wdata,
  input  [63:0] io_cpu_0_regacc_rdata,
  input         io_cpu_0_regacc_busy,
  output        io_cpu_0_inst64,
  output [31:0] io_cpu_0_inst64_raw,
  output        io_cpu_0_inst64_nowait,
  input         io_cpu_0_inst64_ready,
  output        io_cpu_0_inst64_flush,
  input         io_cpu_0_inst64_busy,
  input         io_cpu_1_inited,
  input  [1:0]  io_cpu_1_priv,
  output        io_cpu_1_ext_itr,
  output        io_cpu_1_stop_fetch,
  output        io_cpu_1_regacc_rd,
  output        io_cpu_1_regacc_wt,
  output [4:0]  io_cpu_1_regacc_idx,
  output [63:0] io_cpu_1_regacc_wdata,
  input  [63:0] io_cpu_1_regacc_rdata,
  input         io_cpu_1_regacc_busy,
  output        io_cpu_1_inst64,
  output [31:0] io_cpu_1_inst64_raw,
  output        io_cpu_1_inst64_nowait,
  input         io_cpu_1_inst64_ready,
  output        io_cpu_1_inst64_flush,
  input         io_cpu_1_inst64_busy,
  input         io_cpu_2_inited,
  input  [1:0]  io_cpu_2_priv,
  output        io_cpu_2_ext_itr,
  output        io_cpu_2_stop_fetch,
  output        io_cpu_2_regacc_rd,
  output        io_cpu_2_regacc_wt,
  output [4:0]  io_cpu_2_regacc_idx,
  output [63:0] io_cpu_2_regacc_wdata,
  input  [63:0] io_cpu_2_regacc_rdata,
  input         io_cpu_2_regacc_busy,
  output        io_cpu_2_inst64,
  output [31:0] io_cpu_2_inst64_raw,
  output        io_cpu_2_inst64_nowait,
  input         io_cpu_2_inst64_ready,
  output        io_cpu_2_inst64_flush,
  input         io_cpu_2_inst64_busy,
  input         io_cpu_3_inited,
  input  [1:0]  io_cpu_3_priv,
  output        io_cpu_3_ext_itr,
  output        io_cpu_3_stop_fetch,
  output        io_cpu_3_regacc_rd,
  output        io_cpu_3_regacc_wt,
  output [4:0]  io_cpu_3_regacc_idx,
  output [63:0] io_cpu_3_regacc_wdata,
  input  [63:0] io_cpu_3_regacc_rdata,
  input         io_cpu_3_regacc_busy,
  output        io_cpu_3_inst64,
  output [31:0] io_cpu_3_inst64_raw,
  output        io_cpu_3_inst64_nowait,
  input         io_cpu_3_inst64_ready,
  output        io_cpu_3_inst64_flush,
  input         io_cpu_3_inst64_busy,
  output        io_txd,
  input         io_rxd,
  output [7:0]  io_dbg_sta,
  output [7:0]  io_state,
  output [7:0]  io_cpu_state,
  output [7:0]  io_opcode,
  output [7:0]  io_rx_data,
  output [15:0] io_rx_buf,
  output [1:0]  io_rx_in,
  output [7:0]  io_rx_queue_in,
  output [7:0]  io_uart_buf
);
  wire  ctrl_clock; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_reset; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_inited; // @[NulCtrlMP.scala 986:22]
  wire [1:0] ctrl_io_cpu_0_priv; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_ext_itr; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_stop_fetch; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_regacc_rd; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_regacc_wt; // @[NulCtrlMP.scala 986:22]
  wire [4:0] ctrl_io_cpu_0_regacc_idx; // @[NulCtrlMP.scala 986:22]
  wire [63:0] ctrl_io_cpu_0_regacc_wdata; // @[NulCtrlMP.scala 986:22]
  wire [63:0] ctrl_io_cpu_0_regacc_rdata; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_regacc_busy; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_inst64; // @[NulCtrlMP.scala 986:22]
  wire [31:0] ctrl_io_cpu_0_inst64_raw; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_inst64_nowait; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_inst64_ready; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_inst64_flush; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_0_inst64_busy; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_inited; // @[NulCtrlMP.scala 986:22]
  wire [1:0] ctrl_io_cpu_1_priv; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_ext_itr; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_stop_fetch; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_regacc_rd; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_regacc_wt; // @[NulCtrlMP.scala 986:22]
  wire [4:0] ctrl_io_cpu_1_regacc_idx; // @[NulCtrlMP.scala 986:22]
  wire [63:0] ctrl_io_cpu_1_regacc_wdata; // @[NulCtrlMP.scala 986:22]
  wire [63:0] ctrl_io_cpu_1_regacc_rdata; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_regacc_busy; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_inst64; // @[NulCtrlMP.scala 986:22]
  wire [31:0] ctrl_io_cpu_1_inst64_raw; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_inst64_nowait; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_inst64_ready; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_inst64_flush; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_1_inst64_busy; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_inited; // @[NulCtrlMP.scala 986:22]
  wire [1:0] ctrl_io_cpu_2_priv; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_ext_itr; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_stop_fetch; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_regacc_rd; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_regacc_wt; // @[NulCtrlMP.scala 986:22]
  wire [4:0] ctrl_io_cpu_2_regacc_idx; // @[NulCtrlMP.scala 986:22]
  wire [63:0] ctrl_io_cpu_2_regacc_wdata; // @[NulCtrlMP.scala 986:22]
  wire [63:0] ctrl_io_cpu_2_regacc_rdata; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_regacc_busy; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_inst64; // @[NulCtrlMP.scala 986:22]
  wire [31:0] ctrl_io_cpu_2_inst64_raw; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_inst64_nowait; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_inst64_ready; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_inst64_flush; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_2_inst64_busy; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_inited; // @[NulCtrlMP.scala 986:22]
  wire [1:0] ctrl_io_cpu_3_priv; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_ext_itr; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_stop_fetch; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_regacc_rd; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_regacc_wt; // @[NulCtrlMP.scala 986:22]
  wire [4:0] ctrl_io_cpu_3_regacc_idx; // @[NulCtrlMP.scala 986:22]
  wire [63:0] ctrl_io_cpu_3_regacc_wdata; // @[NulCtrlMP.scala 986:22]
  wire [63:0] ctrl_io_cpu_3_regacc_rdata; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_regacc_busy; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_inst64; // @[NulCtrlMP.scala 986:22]
  wire [31:0] ctrl_io_cpu_3_inst64_raw; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_inst64_nowait; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_inst64_ready; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_inst64_flush; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_cpu_3_inst64_busy; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_tx_ready; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_tx_valid; // @[NulCtrlMP.scala 986:22]
  wire [7:0] ctrl_io_tx_bits; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_rx_ready; // @[NulCtrlMP.scala 986:22]
  wire  ctrl_io_rx_valid; // @[NulCtrlMP.scala 986:22]
  wire [7:0] ctrl_io_rx_bits; // @[NulCtrlMP.scala 986:22]
  wire [7:0] ctrl_io_dbg_sta; // @[NulCtrlMP.scala 986:22]
  wire [7:0] ctrl_io_state; // @[NulCtrlMP.scala 986:22]
  wire [7:0] ctrl_io_cpu_state; // @[NulCtrlMP.scala 986:22]
  wire [7:0] ctrl_io_opcode; // @[NulCtrlMP.scala 986:22]
  wire [7:0] ctrl_io_rx_data; // @[NulCtrlMP.scala 986:22]
  wire [63:0] ctrl_io_buildTime; // @[NulCtrlMP.scala 986:22]
  wire [7:0] ctrl_io_uart_buf; // @[NulCtrlMP.scala 986:22]
  wire  tx_clock; // @[NulCtrlMP.scala 987:20]
  wire  tx_reset; // @[NulCtrlMP.scala 987:20]
  wire  tx_io_txd; // @[NulCtrlMP.scala 987:20]
  wire  tx_io_channel_ready; // @[NulCtrlMP.scala 987:20]
  wire  tx_io_channel_valid; // @[NulCtrlMP.scala 987:20]
  wire [7:0] tx_io_channel_bits; // @[NulCtrlMP.scala 987:20]
  wire  rx_clock; // @[NulCtrlMP.scala 988:20]
  wire  rx_reset; // @[NulCtrlMP.scala 988:20]
  wire  rx_io_rxd; // @[NulCtrlMP.scala 988:20]
  wire  rx_io_channel_ready; // @[NulCtrlMP.scala 988:20]
  wire  rx_io_channel_valid; // @[NulCtrlMP.scala 988:20]
  wire [7:0] rx_io_channel_bits; // @[NulCtrlMP.scala 988:20]
  wire  rxbuffer_clock; // @[NulCtrlMP.scala 989:26]
  wire  rxbuffer_reset; // @[NulCtrlMP.scala 989:26]
  wire  rxbuffer_io_enq_ready; // @[NulCtrlMP.scala 989:26]
  wire  rxbuffer_io_enq_valid; // @[NulCtrlMP.scala 989:26]
  wire [7:0] rxbuffer_io_enq_bits; // @[NulCtrlMP.scala 989:26]
  wire  rxbuffer_io_deq_ready; // @[NulCtrlMP.scala 989:26]
  wire  rxbuffer_io_deq_valid; // @[NulCtrlMP.scala 989:26]
  wire [7:0] rxbuffer_io_deq_bits; // @[NulCtrlMP.scala 989:26]
  wire [9:0] rxbuffer_io_count; // @[NulCtrlMP.scala 989:26]
  wire  txbuffer_clock; // @[NulCtrlMP.scala 990:26]
  wire  txbuffer_reset; // @[NulCtrlMP.scala 990:26]
  wire  txbuffer_io_enq_ready; // @[NulCtrlMP.scala 990:26]
  wire  txbuffer_io_enq_valid; // @[NulCtrlMP.scala 990:26]
  wire [7:0] txbuffer_io_enq_bits; // @[NulCtrlMP.scala 990:26]
  wire  txbuffer_io_deq_ready; // @[NulCtrlMP.scala 990:26]
  wire  txbuffer_io_deq_valid; // @[NulCtrlMP.scala 990:26]
  wire [7:0] txbuffer_io_deq_bits; // @[NulCtrlMP.scala 990:26]
  wire  _io_rx_in_T = ~io_rxd; // @[NulCtrlMP.scala 998:21]
  NulCPUCtrlMP ctrl ( // @[NulCtrlMP.scala 986:22]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_cpu_0_inited(ctrl_io_cpu_0_inited),
    .io_cpu_0_priv(ctrl_io_cpu_0_priv),
    .io_cpu_0_ext_itr(ctrl_io_cpu_0_ext_itr),
    .io_cpu_0_stop_fetch(ctrl_io_cpu_0_stop_fetch),
    .io_cpu_0_regacc_rd(ctrl_io_cpu_0_regacc_rd),
    .io_cpu_0_regacc_wt(ctrl_io_cpu_0_regacc_wt),
    .io_cpu_0_regacc_idx(ctrl_io_cpu_0_regacc_idx),
    .io_cpu_0_regacc_wdata(ctrl_io_cpu_0_regacc_wdata),
    .io_cpu_0_regacc_rdata(ctrl_io_cpu_0_regacc_rdata),
    .io_cpu_0_regacc_busy(ctrl_io_cpu_0_regacc_busy),
    .io_cpu_0_inst64(ctrl_io_cpu_0_inst64),
    .io_cpu_0_inst64_raw(ctrl_io_cpu_0_inst64_raw),
    .io_cpu_0_inst64_nowait(ctrl_io_cpu_0_inst64_nowait),
    .io_cpu_0_inst64_ready(ctrl_io_cpu_0_inst64_ready),
    .io_cpu_0_inst64_flush(ctrl_io_cpu_0_inst64_flush),
    .io_cpu_0_inst64_busy(ctrl_io_cpu_0_inst64_busy),
    .io_cpu_1_inited(ctrl_io_cpu_1_inited),
    .io_cpu_1_priv(ctrl_io_cpu_1_priv),
    .io_cpu_1_ext_itr(ctrl_io_cpu_1_ext_itr),
    .io_cpu_1_stop_fetch(ctrl_io_cpu_1_stop_fetch),
    .io_cpu_1_regacc_rd(ctrl_io_cpu_1_regacc_rd),
    .io_cpu_1_regacc_wt(ctrl_io_cpu_1_regacc_wt),
    .io_cpu_1_regacc_idx(ctrl_io_cpu_1_regacc_idx),
    .io_cpu_1_regacc_wdata(ctrl_io_cpu_1_regacc_wdata),
    .io_cpu_1_regacc_rdata(ctrl_io_cpu_1_regacc_rdata),
    .io_cpu_1_regacc_busy(ctrl_io_cpu_1_regacc_busy),
    .io_cpu_1_inst64(ctrl_io_cpu_1_inst64),
    .io_cpu_1_inst64_raw(ctrl_io_cpu_1_inst64_raw),
    .io_cpu_1_inst64_nowait(ctrl_io_cpu_1_inst64_nowait),
    .io_cpu_1_inst64_ready(ctrl_io_cpu_1_inst64_ready),
    .io_cpu_1_inst64_flush(ctrl_io_cpu_1_inst64_flush),
    .io_cpu_1_inst64_busy(ctrl_io_cpu_1_inst64_busy),
    .io_cpu_2_inited(ctrl_io_cpu_2_inited),
    .io_cpu_2_priv(ctrl_io_cpu_2_priv),
    .io_cpu_2_ext_itr(ctrl_io_cpu_2_ext_itr),
    .io_cpu_2_stop_fetch(ctrl_io_cpu_2_stop_fetch),
    .io_cpu_2_regacc_rd(ctrl_io_cpu_2_regacc_rd),
    .io_cpu_2_regacc_wt(ctrl_io_cpu_2_regacc_wt),
    .io_cpu_2_regacc_idx(ctrl_io_cpu_2_regacc_idx),
    .io_cpu_2_regacc_wdata(ctrl_io_cpu_2_regacc_wdata),
    .io_cpu_2_regacc_rdata(ctrl_io_cpu_2_regacc_rdata),
    .io_cpu_2_regacc_busy(ctrl_io_cpu_2_regacc_busy),
    .io_cpu_2_inst64(ctrl_io_cpu_2_inst64),
    .io_cpu_2_inst64_raw(ctrl_io_cpu_2_inst64_raw),
    .io_cpu_2_inst64_nowait(ctrl_io_cpu_2_inst64_nowait),
    .io_cpu_2_inst64_ready(ctrl_io_cpu_2_inst64_ready),
    .io_cpu_2_inst64_flush(ctrl_io_cpu_2_inst64_flush),
    .io_cpu_2_inst64_busy(ctrl_io_cpu_2_inst64_busy),
    .io_cpu_3_inited(ctrl_io_cpu_3_inited),
    .io_cpu_3_priv(ctrl_io_cpu_3_priv),
    .io_cpu_3_ext_itr(ctrl_io_cpu_3_ext_itr),
    .io_cpu_3_stop_fetch(ctrl_io_cpu_3_stop_fetch),
    .io_cpu_3_regacc_rd(ctrl_io_cpu_3_regacc_rd),
    .io_cpu_3_regacc_wt(ctrl_io_cpu_3_regacc_wt),
    .io_cpu_3_regacc_idx(ctrl_io_cpu_3_regacc_idx),
    .io_cpu_3_regacc_wdata(ctrl_io_cpu_3_regacc_wdata),
    .io_cpu_3_regacc_rdata(ctrl_io_cpu_3_regacc_rdata),
    .io_cpu_3_regacc_busy(ctrl_io_cpu_3_regacc_busy),
    .io_cpu_3_inst64(ctrl_io_cpu_3_inst64),
    .io_cpu_3_inst64_raw(ctrl_io_cpu_3_inst64_raw),
    .io_cpu_3_inst64_nowait(ctrl_io_cpu_3_inst64_nowait),
    .io_cpu_3_inst64_ready(ctrl_io_cpu_3_inst64_ready),
    .io_cpu_3_inst64_flush(ctrl_io_cpu_3_inst64_flush),
    .io_cpu_3_inst64_busy(ctrl_io_cpu_3_inst64_busy),
    .io_tx_ready(ctrl_io_tx_ready),
    .io_tx_valid(ctrl_io_tx_valid),
    .io_tx_bits(ctrl_io_tx_bits),
    .io_rx_ready(ctrl_io_rx_ready),
    .io_rx_valid(ctrl_io_rx_valid),
    .io_rx_bits(ctrl_io_rx_bits),
    .io_dbg_sta(ctrl_io_dbg_sta),
    .io_state(ctrl_io_state),
    .io_cpu_state(ctrl_io_cpu_state),
    .io_opcode(ctrl_io_opcode),
    .io_rx_data(ctrl_io_rx_data),
    .io_buildTime(ctrl_io_buildTime),
    .io_uart_buf(ctrl_io_uart_buf)
  );
  Tx tx ( // @[NulCtrlMP.scala 987:20]
    .clock(tx_clock),
    .reset(tx_reset),
    .io_txd(tx_io_txd),
    .io_channel_ready(tx_io_channel_ready),
    .io_channel_valid(tx_io_channel_valid),
    .io_channel_bits(tx_io_channel_bits)
  );
  Rx rx ( // @[NulCtrlMP.scala 988:20]
    .clock(rx_clock),
    .reset(rx_reset),
    .io_rxd(rx_io_rxd),
    .io_channel_ready(rx_io_channel_ready),
    .io_channel_valid(rx_io_channel_valid),
    .io_channel_bits(rx_io_channel_bits)
  );
  Queue_1 rxbuffer ( // @[NulCtrlMP.scala 989:26]
    .clock(rxbuffer_clock),
    .reset(rxbuffer_reset),
    .io_enq_ready(rxbuffer_io_enq_ready),
    .io_enq_valid(rxbuffer_io_enq_valid),
    .io_enq_bits(rxbuffer_io_enq_bits),
    .io_deq_ready(rxbuffer_io_deq_ready),
    .io_deq_valid(rxbuffer_io_deq_valid),
    .io_deq_bits(rxbuffer_io_deq_bits),
    .io_count(rxbuffer_io_count)
  );
  Queue_2 txbuffer ( // @[NulCtrlMP.scala 990:26]
    .clock(txbuffer_clock),
    .reset(txbuffer_reset),
    .io_enq_ready(txbuffer_io_enq_ready),
    .io_enq_valid(txbuffer_io_enq_valid),
    .io_enq_bits(txbuffer_io_enq_bits),
    .io_deq_ready(txbuffer_io_deq_ready),
    .io_deq_valid(txbuffer_io_deq_valid),
    .io_deq_bits(txbuffer_io_deq_bits)
  );
  assign io_cpu_0_ext_itr = ctrl_io_cpu_0_ext_itr; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_0_stop_fetch = ctrl_io_cpu_0_stop_fetch; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_0_regacc_rd = ctrl_io_cpu_0_regacc_rd; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_0_regacc_wt = ctrl_io_cpu_0_regacc_wt; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_0_regacc_idx = ctrl_io_cpu_0_regacc_idx; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_0_regacc_wdata = ctrl_io_cpu_0_regacc_wdata; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_0_inst64 = ctrl_io_cpu_0_inst64; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_0_inst64_raw = ctrl_io_cpu_0_inst64_raw; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_0_inst64_nowait = ctrl_io_cpu_0_inst64_nowait; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_0_inst64_flush = ctrl_io_cpu_0_inst64_flush; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_ext_itr = ctrl_io_cpu_1_ext_itr; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_stop_fetch = ctrl_io_cpu_1_stop_fetch; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_regacc_rd = ctrl_io_cpu_1_regacc_rd; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_regacc_wt = ctrl_io_cpu_1_regacc_wt; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_regacc_idx = ctrl_io_cpu_1_regacc_idx; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_regacc_wdata = ctrl_io_cpu_1_regacc_wdata; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_inst64 = ctrl_io_cpu_1_inst64; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_inst64_raw = ctrl_io_cpu_1_inst64_raw; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_inst64_nowait = ctrl_io_cpu_1_inst64_nowait; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_1_inst64_flush = ctrl_io_cpu_1_inst64_flush; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_ext_itr = ctrl_io_cpu_2_ext_itr; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_stop_fetch = ctrl_io_cpu_2_stop_fetch; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_regacc_rd = ctrl_io_cpu_2_regacc_rd; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_regacc_wt = ctrl_io_cpu_2_regacc_wt; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_regacc_idx = ctrl_io_cpu_2_regacc_idx; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_regacc_wdata = ctrl_io_cpu_2_regacc_wdata; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_inst64 = ctrl_io_cpu_2_inst64; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_inst64_raw = ctrl_io_cpu_2_inst64_raw; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_inst64_nowait = ctrl_io_cpu_2_inst64_nowait; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_2_inst64_flush = ctrl_io_cpu_2_inst64_flush; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_ext_itr = ctrl_io_cpu_3_ext_itr; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_stop_fetch = ctrl_io_cpu_3_stop_fetch; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_regacc_rd = ctrl_io_cpu_3_regacc_rd; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_regacc_wt = ctrl_io_cpu_3_regacc_wt; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_regacc_idx = ctrl_io_cpu_3_regacc_idx; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_regacc_wdata = ctrl_io_cpu_3_regacc_wdata; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_inst64 = ctrl_io_cpu_3_inst64; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_inst64_raw = ctrl_io_cpu_3_inst64_raw; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_inst64_nowait = ctrl_io_cpu_3_inst64_nowait; // @[NulCtrlMP.scala 1003:12]
  assign io_cpu_3_inst64_flush = ctrl_io_cpu_3_inst64_flush; // @[NulCtrlMP.scala 1003:12]
  assign io_txd = tx_io_txd; // @[NulCtrlMP.scala 1004:12]
  assign io_dbg_sta = ctrl_io_dbg_sta; // @[NulCtrlMP.scala 992:16]
  assign io_state = ctrl_io_state; // @[NulCtrlMP.scala 993:14]
  assign io_cpu_state = ctrl_io_cpu_state; // @[NulCtrlMP.scala 994:18]
  assign io_opcode = ctrl_io_opcode; // @[NulCtrlMP.scala 995:15]
  assign io_rx_data = ctrl_io_rx_data; // @[NulCtrlMP.scala 996:16]
  assign io_rx_buf = {{6'd0}, rxbuffer_io_count}; // @[NulCtrlMP.scala 997:15]
  assign io_rx_in = {_io_rx_in_T,rx_io_rxd}; // @[Cat.scala 31:58]
  assign io_rx_queue_in = rxbuffer_io_enq_bits; // @[NulCtrlMP.scala 999:20]
  assign io_uart_buf = ctrl_io_uart_buf; // @[NulCtrlMP.scala 1000:17]
  assign ctrl_clock = clock;
  assign ctrl_reset = reset;
  assign ctrl_io_cpu_0_inited = io_cpu_0_inited; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_0_priv = io_cpu_0_priv; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_0_regacc_rdata = io_cpu_0_regacc_rdata; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_0_regacc_busy = io_cpu_0_regacc_busy; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_0_inst64_ready = io_cpu_0_inst64_ready; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_0_inst64_busy = io_cpu_0_inst64_busy; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_1_inited = io_cpu_1_inited; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_1_priv = io_cpu_1_priv; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_1_regacc_rdata = io_cpu_1_regacc_rdata; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_1_regacc_busy = io_cpu_1_regacc_busy; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_1_inst64_ready = io_cpu_1_inst64_ready; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_1_inst64_busy = io_cpu_1_inst64_busy; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_2_inited = io_cpu_2_inited; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_2_priv = io_cpu_2_priv; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_2_regacc_rdata = io_cpu_2_regacc_rdata; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_2_regacc_busy = io_cpu_2_regacc_busy; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_2_inst64_ready = io_cpu_2_inst64_ready; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_2_inst64_busy = io_cpu_2_inst64_busy; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_3_inited = io_cpu_3_inited; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_3_priv = io_cpu_3_priv; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_3_regacc_rdata = io_cpu_3_regacc_rdata; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_3_regacc_busy = io_cpu_3_regacc_busy; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_3_inst64_ready = io_cpu_3_inst64_ready; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_cpu_3_inst64_busy = io_cpu_3_inst64_busy; // @[NulCtrlMP.scala 1003:12]
  assign ctrl_io_tx_ready = txbuffer_io_enq_ready; // @[NulCtrlMP.scala 1006:16]
  assign ctrl_io_rx_valid = rxbuffer_io_deq_valid; // @[NulCtrlMP.scala 1007:16]
  assign ctrl_io_rx_bits = rxbuffer_io_deq_bits; // @[NulCtrlMP.scala 1007:16]
  assign tx_clock = clock;
  assign tx_reset = reset;
  assign tx_io_channel_valid = txbuffer_io_deq_valid; // @[NulCtrlMP.scala 1009:21]
  assign tx_io_channel_bits = txbuffer_io_deq_bits; // @[NulCtrlMP.scala 1009:21]
  assign rx_clock = clock;
  assign rx_reset = reset;
  assign rx_io_rxd = io_rxd; // @[NulCtrlMP.scala 1005:15]
  assign rx_io_channel_ready = rxbuffer_io_enq_ready; // @[NulCtrlMP.scala 1008:21]
  assign rxbuffer_clock = clock;
  assign rxbuffer_reset = reset;
  assign rxbuffer_io_enq_valid = rx_io_channel_valid; // @[NulCtrlMP.scala 1008:21]
  assign rxbuffer_io_enq_bits = rx_io_channel_bits; // @[NulCtrlMP.scala 1008:21]
  assign rxbuffer_io_deq_ready = ctrl_io_rx_ready; // @[NulCtrlMP.scala 1007:16]
  assign txbuffer_clock = clock;
  assign txbuffer_reset = reset;
  assign txbuffer_io_enq_valid = ctrl_io_tx_valid; // @[NulCtrlMP.scala 1006:16]
  assign txbuffer_io_enq_bits = ctrl_io_tx_bits; // @[NulCtrlMP.scala 1006:16]
  assign txbuffer_io_deq_ready = tx_io_channel_ready; // @[NulCtrlMP.scala 1009:21]
endmodule
